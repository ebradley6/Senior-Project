��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z��4֬��9�A��;Un��Gh[�����<�#�L�-8�o����X0v�c�4��S�`U��� ik�{=�g]�C�+a
>kN}%]q�]���g��k���Y1b	 ���5��G��r>��T�CF�h��PNdi��NS�rd�j�FN��!X�fɅ=&t]������0��R��1�b"�܍��#��LJC�G��o�à���zz��c��Iq#����s�h��wb�¯(�"Iɇ�օw¶}��s�n���^�AI��������`B *?z�/��Z�/�bp4�-�~�L����>ҥ�x�&kD���F"py��B���ͪ�*1�@�}��*�W�q̄��9��[XC�{\['{�w��$�d�$L���d�t��S��"	x���mե��9*��:��pT�<�:꾖����ҌL�q@�-�=��
��\3�&�ϩ����|@�������c$�m�@KaY�Ҙu;�An�UNh����Z��o7���������l���sK���> 3߀�:K����D���ޭ?�	��t�\s�O��(�މw���#������N��QE:l�^��R[o�܀Ms�����u�§S?�F�����#����JE���=�b5�A-�:ʚn%������}mE����|��K�r�r
��~e��k6x-C������؋B�� d@yb�m�_.�o��,"�V{&����tI�
`�����U�?�tI�)��\M
l�.����Z�M�u"v�(���;|�#L�7����s�o���O�^oRY�Y� z����S�׫�D͚t����|�χ�y�*����B;�~�v׃h����21�o�k4��&Aߠ9&�~��a$�m1t� ʄ�a~ր#J.���k��(���A�<q�� ER��ٚ�&��&�&/����3������+�@��c/�_]Ds��������`�*�?�t����y�"��g�?A)~��tt�t��.ed�d1���ȑ��ʼ�Xp\�Bs����[��})��{&�RY=4U�U�,�F�ךд�o�m3��߇`������c�HS�����嶌�.�_KSU"�W�Z
S;�6h�V����n7����{Ӯ;�[��4��^Q�.w��O�c���X�)(�n�Ù��kG0J��=Ȼ4�G�BcD�K��A�"Y/l���H�x~{e&8���"Ч>\B�t�6:y�%U���u��͇�8��s^��\ҩQ��J���U�f��G|Eg��lZJ\�j����q2�.�6���(t����ɗ��WN��#�-%���^X/ۍp�����i�ӝ���PnC�(�����Ԕ��{����h�b��]�7?���Z�H�QyX���})�cbXљ��=}!Z�c]�ӡ"��{����0�y�B3F��~3�lI3cLͱ H�I�x\E�&�/iVciR��ſ���A��a��%���o�F?���W�bѼKn'Y*SM�o���)Y��s�Ӆ��9f1����;)d@EA>��H��5|'4~�
z����6�n��
�w�%�!����n�!�=;CK/
�A�л>�ê�tt�`� �Z͠X3i&hY�-��zem�Dy�#E��g��G�߁���)z'������AO�D�aP�����{<��<�K��:{_��ٗ��;��;�e�6	�u���mZ��e��� G`��_4t���)Z{uw�~�D�i<M�ܵ��[vĔ�k��v��f��������A~�<�JS�o�cM��"�G ��e�+�[=�?1�2I�H��R��%s��w��Ȩ�#�][���Ts����̎u�b�s�����g�te��>�ޖ�z�� Z�'y��1"3zz�#[7�aI�g�Q��#Ũ���G@M�����2��./P>�f@��'�C���3:�l�V@��ťd�4J�UP�#�Qi��n���m��>�i>�d袴�,�&ݦ�c�I;o�Q&5�|�G����� 3}S"���a	~�Э$�+F�N�L�����T=�?w�x��v>�VU��FO��|�����B^(�xu��V3}�"N�7k��b�3�v~����A�c��+��j������#[�ue�D���J�_'�߱k4��!��D{�nd��?�<	���KD^R�ud�X��en1���S`�G�G��F$��%�J�W/�nA�H����K�$Q��H*NR�I�����Ǯ��zy+y�)(�(���@a�q���.)N#�(0��?d���p'H�B�i�}�#}���.E�#C�>�����:ϹNS�8������QGl���� >|�M��8�T��0�K��rqA_v�[�{ń岰T>*�q�澏2���h�s
���d*Ym��y��:�\K�E�Ej� ��`�Q�;>h�f��i8�
=�"�:�ov-������(*��}O�j�}� �$jV/��>�Ky������r�ei�X�j �0�4�~�{��~j&�nk2����e3D�T:
����#�ͥ::ZzJȉtɖ�}�	ܴɰ�"|ؗ�9�K����H�Ҋ6z~%�X��`���jj}M��,���)h*�e�wEtb�~p�*�fU�NTt���A��宐�F��D
��_��l��X*.�+f\�AK��#s���L�F�@��Q)~��b���J1�4���x|2C�:��R�1�_�b�!��#T K��r(��W��4?jtX�ep���!��wW.�������6v��rPEy@aQ6L���*֣yF3�x�O�O��S�;]�cxj��A�{�^�W�ʅ��m�6�-&���I����d���;��?nU����o$[��c�v&d-�W*�K	fB� ���/ ��,.C�k�+���1��W��}R u���c����R�7�Pg�b$�w�8j%�;!��DܦT@��_�~��(��T�o�A��F�t���F��K���܃��s��GL8�ئ�2=T�K ja�?�G���Tn#'�G�����Ԛ_=\�Ҧ��bb>�+�}�L�o�?<6���]������� AT>8���\?�ck�3�7)V���4�q�q	��Vr}�*��N����+P���4~X�5�h��.�o��J����$IkBW�Au�[����s\3)c}�d��$����wT�q�z��O}�f�\+������8�$7�cQ�<�g���h!��"]���k�41��sC�����X��ΰ����,�My��ē>�����Z�2��J��9χ�E�8l�^(��b�����3�@Ê1�4"Qh�e4~<��?0/��Ǎ|�o��/Ĵ���+
hl;!�(����+FxIR������=�~��y~٤�̱K�!>]�.�0,�^KR��u_�S	��d��~�+cXg�����9aYK��һ��g('GHg�̟V%/���M���'�M��*\��G�ת)��؇Pa|�L7��,�fO�q��{�
�$|��ұV<��QAW	�!:C)PF�c�9�e)@�UagP3kh�^`�Ͷ\y�2�j�qo���ggBs��	���㫱kϏQ�q:\�F�R�F� /�l� �(������������F2��\J�y<쭲��G��J�CYş����#����;�Xg���~�SF��R��&Tn��O+�^3�Q��� "b��D�1ef��y�.����vt�r�ؗ�M��Wҹ��fs�!�;�B�nIk��6� n�re�$�'FL�>�P^䘥%�oN�`����1rlb�� �K�셪�IW���|SI�%�bu1/0�,�n~�
&��?�A�%o�.h0��bO�1����*�?�ZO�v>��c��z��2$�@����2#�/% .���x/E0��+�[L�縚��y�qH����yL�uT
c�U47(	S�Oj��b�n����X��8ڿ�-��>���v�п�;hK�f΂����j~��Ѝ��N�R���V�?���K�N�f4�/A�p��g�*YW@���Z�m������3��2x�f��39*�BqX��3���D����_�����6��p�%)�­���d�!]⭬b��ݐ8kZ�G#J^�_�Z�&L/���pc6�Z'^�{�o��*)�� ־l|�մ(JS1���̼�)�|'ۖ�	W�F-.�y
�Q'0�(�����f���?_�0�|�4O^���8�{��L�P�C��=��2�OZ�NM�%MG͐�N��	Lɳ��^0G���m�B�����MQ�)�4���}����8y0��5�,������\�����wN��^ ��p�)���g$ ^��a�?�q@��y�-��w�;P���$�cQ�3����o�.y��1��M[ Q{�k��x�Yc���/�c�y�����r�pw�,�f���} [xo�P�tn�<��
�M�k�_�?�����nO��-��g�A�$>��tHJ��8非�~{2���1/`�:�y�2�_��.n�~��L\�Ix����L	x�a��q]�6��i�|��PҔъ�]��������J]$}�]{���ա;��;���=� �~�t�-���T�M-f�,���������}f�Ü���s~��6g�
����^��a��_h�~\�38?��namEX��-���T��ҷ�8|+t���o]�v{�r��R�W�:�S�
��.��@-8 g�� �E��Sf�V|���#�o\c��]L���ߠ����(
�]5����w�h��_���9��UH'RQ���"|�����j!�n��1W�[Ir�V�����=b�XmLQ�z�C������x`u����x�z
\�>�W�{�W�.$�RE�O���/cՄ� �ph�u4���ٺ,s%�I`��!��� ��Z���1���9���şԸ�)�/�Q��m��*Z����7J�b̃F%[�镨�H�4L�5r~��"a�ɢ��;z��S��-�_?��{o���� xA��v6�pP	ѢrZk��+!(@���i�	{�rӠ������~z���q����ZΗ�u���'�.�1���`gk:�|�QaߢL�	�
w6�)����&`������f��T�kfV1��һJv0�b-3T h��C����[�2뭮NM�01ue!�Kٜ45�2 ���v��,6D{�q�h��:�b��
];d\a�Е]%���c��Qc�hz@�o�o%p�2��[�����7�56w�qF�4�^v);�a����j+Yꢢ [D@��.�i䯃���t�mfM$��i���JM�*o!���z�3Ae��1��SiE���j�.�ZC]��ui�E<=g_6�n����>F^��������{����9����/#��իݹ><\�\?��I�A�5*��}p���}h�)X�qS5'��U�]C��Z�^��>ש�c��|�s'����J�!�V���$}^ŧ�,�w%���TzKD�� ��hF"���Ef���d)� �q��b�Һ���\M����+�y:.N|΢�,i�;e2!���g"�Ƚ�\t=�=-������Ey�xv5P������ncއΰ#�a�R�1�G���#Ѕǎ���X'
!ݖ�|�F�%%����t�S���ε�'XG=pL^2)Zon��i�D��2���d|=�v��D@���?������H���P�Y�k��-	򿕍�N���[�*8����,�����7�\�W��ù_V���>�$bt�kO�ڭ��gKC��ڞ���*��� v�0�v������v�䈏2�H	�@�8	�~�󹥤�A[L��|f%l�we<Q4���V��yB:�yW���m|�U"�'�N2��3^�Ε�z���F���u+lW#D
;�C��8Z��e#j��!�Y_ϯ�R+�lY(��n��nu��I]�^��Ӣ��a5�@�����.���NTޝ�;F:I��B���n�����h�
B҄�R�t%������I�Yi�� 4��v�B��'��)��I��唵4��*��n`{E�4Q�� ��^���-�L���d07]uOe��R1��w2���@�-�Q����a{N�щ�7���]Rq-P:�Z+z-`�H���xC��n2k/�����R}B����O4�]�ŸypeQM?@c������o':�Y,o螰�%{�PY�Y�5�Gֱ����1�B��f}��-p�C���@]|���f�l��Qij��.���LiR�WW����4�.̑�`�g'N�<�&֙�}�i�`!����x�L�� ח�Z����<y������;�Zz�v[i٥_a�n����xLN �Qm@i����*Jϰ���4�����?�ze�d�?���s����&M�Z( ��e�-g0��y�@�5ߵS%�%Qe�B����$�k����AH�i��!(�r����7��Kgx�~���3cϋ�k��L��4��x����&��u
pi�BVn��n�_V�����D�sSt�i���K�h�`�,�I�Or�ehb�(�.�3ѥCf������+�y5�T�E�?TX�*F�V�}a˷_�v~���������<�:TP�'-�'R��AD���9�R���g���Nj/O���C4��Ʊ@�J�[b#��=�8v���-��$ML�����S	���]H�_�m���c�{Ԇ(���O|I��g�´R��#��lOz��0A7��M�q*ĭ$;��^��V�+���-w�Nk-���H-Z5��R�������8��)��~��,뚻*uœ��`�d�/[#���6�?�`��14@�%dα�b�5nʜ��ĸvi��!���w�*�<�����7�1w'���2�b��t�3g���)�s���A�r��2$�)�-2�G!�J�ɼ������&�}:T����a2��a!�����Z�m*��O�;���u�	����ǗT�������Xx�E{7�������p6O��x������O��+K����^ �:`r|9����j��s
}��瞝�K3A�
�˧@���)��z���"���XM)�(!A�����9��,�+�	.{�U�sz��0S��/ŪTjP^dzygZ}x�s�p7�]�4��d߫���D˴d�ȔZ���>d���?ŕ�,��Ƽ9v��j����5�#[�zA���fV���
�"T�~���f]p֩����|2���c�FB��l��0G����QoY��B�>����N.)ʶc~C�7V�P�_2���6�I74���6�E%ȵ��,����=']%rze7W�Vܻy��E1��#����2kZ����p�$�&`�o[n���;�}��{���bʠ$� �J8#�S�_�k��	���P�a�OX覯���ߟ�~_����S�{��wt�aU7p�4}�Xo�֚�V �/
�S	�Z8���㖹��'�)��T~�F�+��Ϭi���A3�1���bN��eπ�/������=0�H)�^P`_�Dm�����A��IKRF ���M*]28�d�!�ɛQ�h���i�3�:c��xR�o咯�#5K	Ӓ_��s���z���ꪗ[���!�>�ѣ�?i V/A��y����Z��* B�,ʽB9 ��Or�۲���_���m֍��Q����B�a҅��ÕR�O�>��k�O��j^�`
Z�ݢ�E[�p�^jm./
������s�;���T��-�$ӹ�]��a��{�S��.�[q����XH���<�ʋ��>���p)���o�^�&c��W���Y�Uz�4ŭ\���j���YyÄЂ�IT�ؾ+��6��as�� .�FGz�&rrqey�ռ������(���Zpl�eF.��(�2�/�}P-���Ip�Qo��s=��#��ڣ�;E���ݹ� +�BP��!i#"�A��A��hI�ڞ�u��7�/．\N��ߧ��Q��S�3������-�HK�2�퍸�^�	���oϐx���Ƙ�R����t�Ӽ����9d)����� ܨV��������e$˕�)�t*�����R%OT��.�:�'�7�<V�U�~�2	�W���Ӝ�-���uO�����XQ,���@��c�YJ�M��"0q�t�@?�]��� |�: [2��@:i��ǥ�_�d�_U����`Y�6�d�0D������ƀ��AqG���hr�R���g�Q���n�zr�R=B�E+�$��Ûbs�������㼦��I����^�ׅe���}k�x$�p��D�
p�܅����@�4�W��x�}��:;h�4C�~d��kw�I�)X5�G�������-2��_�"���=��	m��?����RRǻ�<>�5��	u�.�{�}{���pK`��,+�$:�>��F��Jv��Ċ<��ec�%�7{8�+H����!R��;���|8f|%_�qI���s(�o{WJ=��{󉚃^�v'�U��m�U�^xي<���$6P��������%lMV;�o�V��~Y%6�8dታ�A���Y�}3v_��:����Ҿ�h3��t܈��䖣9��b�6=>��zU���n�ȭR��>��a�2��OW0���nT���4z	��P������|���۴��P���m�(�����1 =ť�1�s��������V8����HDW��#q�����-��y���7ɿB>[��i��4�Fy�v~��h�ֈ�m��`�\�`a��v���ok�!_/3����t =v�b	�M�n��s.8K-�Pa0�aL5P�k1P<]'=j����#,�]O/��¶�Q*`QY7�^��ɸd��>�o�-té���׬ʽa!�>m�A�xI���9�b@Vq�v������q��CC�?y�`��[̻@@���s��5O���H������nk;��Ҟ�e;]���밒��XB`��d�ؑ��	�I^̵<j�w0�o	�C��f�!E(���}�4��Qi	>�������u)�̸����rD�d͠�Z �a���s������V<z���v�}τ{���]���劷�]�Ϣy֫u��]������qf���������3p \ͳ��UXJ_v�A�x���x�*�ޮ��~�N8�J�����7e����*-m<�����XO�SM<B 0B6����MBQ���5Ι�1��锏M����zk�i4co7��N֙u��Cp��E5k1Ϧ��M{��O�"I5��W�
��B˓?�K�o]�@0��m�mb�rZ5�C��X�,�����Lq�xHzn�SZ	R)=g�;,�o������̭�eǊ����X�=,�d:�Sm�BIH�\��	��W��繁[������܁�m��Y9p/yC�ٴK���|3G��]]�!��ဥ��Mh	��W~���oq0T��
��Czkfn
���^�*d�@4';DZ�����|��)�}][�UMwf7�(IS�K�i�Bg<��:�dS21�Џ�ڊ����RE�=���D^�`�*'ʆu���z�
��l	�Kƀ��&[e[�9��㕁;��#r�E���^��r?���*���kΩM1���PS���FF�P}�&�}Q�&�W��F��c8�L��>��	�}(-T�b�	.1����7��;�ơ׬%�V�5|vx�1���C��6F:�n;��B�Wq���m� ��C�+���z�`�ec���Gv\:jh��62���, �d~?����,[3b�l���M�����X�̜����	��-`�H�b�e�딡��AS%dI+Q:%�Q��u.�X�i�vv�>�����+��3��${�{t��~��*�g���`/�\<�"�a�֊�����F?����!�_lC+���5\O�@��C��dO�&gf�_�(>��_#�6�r���Ƕ��ۻ�FnV�&G��#�E�����z�`J�e��aRi)�S�^��1��f֑n�p)��T8&���j�]�np^5�*g�K^� H*$tZ1�`
V�F1M�VM�ѩ�Y��{�\G��E�L" ��D�\�6צp�� #X��#̒�^Ig��s��^`��X�\��hxU�W�<��3���Tk��U
Q"G��g�D}�VD���fA�3�8,.N�����헦A�̡��u�_��O`�in��$�y�ڈ�&��Q?��eo�/*n����Q�NJ����_J3�����%X���#�?�xUOS����B{^�i�}5m�M:�igSN��?��6�M*�>�j�I�ã9|��@��4#���_�E�t�.���t�3�N����C� ��|�h ����ܳ R�\��F2w?^�]�H9�Z�b�u6���Ib�ꍓ�V��?M��;�7��k�2�hi�MN ��kT̲�����2(kyi��'@$y�3�\KE��͍2`�{o��
߅��4O|�p��C`]�u�[�AW?�>�z!�G��fsC�W�c1�x���l�n,� j�F�)&L���ݙP��>��Ρ�~��:�ǲ�\�=�d�����u{ͷ.�A�ckr��Ic�o���ҵlZ���;�"�{���AԦP։�-ǘ�m�)���<�����6b]�Y.�1_Ȣ�f��r�:dBW��a����J������pW��0&���/:��������f��{�� n�V��6:�E� ���׶$3i��"�+@Г�t���A��P�����>BK��z�y�P���9�)_ҹ`4d������5��Y��R}��a�Rg���H�*zi-�z{xe[�H��
�����/�3h�!Z�3�[�Qv�to�-S��!�{�+]�����S�����f~R�������HK�>�+��ED��ݟH�v;3�C&�������H��Ņz�&d�/�F�$�	HZ�\��~Uy7��ƻ���j{j,�|i:q^�I7}N��q.����A�N��绨�"s�[����3�MҒw_k!��		C�񿛷���!:D�d�unį�r@��EV�n��7CL릈}�>wC�!jA���� �l)eS�{�����⑪̨�q�/"�H�����H/|�Ȫ��ݼ6[�'�+6���|X�˴I�^D��L��II��~��f<U�~���_"���3�����3\.j�.EϬ�H�R�d�i�;��e�Z�1�t�\J̠_�� �88�#AS̹��T���E"1HW6ͅ����wC1�:U�f����-_�I	ͩr����n7��d+`BN\`ڎ�������H�]���4Co�|݌����Z_Lq3�l��;i���.����^����x���j�V�hCr�����'�<��:�|9Z,�QGH�9��HC���E��S�S�@l�B��y"��	<����n�qg���\O_M@�M}2���tr�4[�M�$�sh��OY�{� �!Y\��kqΚ^呸�6K�\dv��F��B�j�Kdv�$�F���0XM�U/n�;E����W�����1�t.���
_���E'�_I��<�]>�\��T��B��/%#>��?z ��q�,�<�)�o�U
����)�ǿ�h��v�� ��"�_��0O�L�q,6.'y�_2�ʍ�{N�k�
Lr$��G�>�D�`Kd�٤��S�>�n��r1A#� �5�}�l>A`-�u9���_Í�s���*�H��1�1����&����r�5�D�a\��'W�D��GO��-P)�j�~L9� z-�8�a��>>�Y�����t�N��!S���bp��}O̟�	|��N���K�C1���B�C7���'!cd�>�[Do����F���&l���j^���A��u�9���YTB���(4�?i�<몼�"k:MT<$�*7�ChH�rN�Os{EH�5�
���$R�N��pS�ڞ ���ʪM��#�&3L��[�&�����+%oY��C��Kw�}M�\g/	��+��W#'�~�as�vO�4��|���ұ̥Y`�7���(�Rبصd�&�Ox�	�o߶"oU�9��P�0�a>jG���W�Ar�g�`6{bR��=���|�ίC���EK���#['���'����y�*I5��}���ɯ|/�X�Oc�*��B��L�Wy��p�����x�[@1�)�e����J�`�Om�����}A0���/=�Cs�`�؀t�"V^�(�~Gz����������O�N���3Զ�H|�8�+\]^���8�bN�����;�1�ms(�GK4��m�wc��'ݺ��B�@rd븠�KE���$��;���3EC�x���YT�j!��Չd.jZ��]l(����G�M�ag��{'S���T�6��=�m��fe���9�<��3F�� �)��&��6�%�G��[���υV=��7@o���\y�d�$b=��j,b��۷���w��I%ud(�Χ�C8�8.����)��Uqx!˘�~Ȳ��S�7ȧ��E	$�*HbJ�|�Ӵ��>e�0׺���y3e��-:e��`=rFk�� ���(d�HM_��1HS��[����0�sFD?y⃳;�+'	�C�,*$���[E�Z����"��E����Nv���\,������
�te��o�{�@������7>+��pM�?���W4�6�@�z��-o̊>?@���. C%P�I��月De��褎)䕸��a;����3p�5���� �̘Bw������p�* �V~Ҏ�d��"��C���+A���?�W���~�q���/����	;B�����ECgī=�d����E��켶L��so��&�<@%j�"ɂ�LH���ՅC@w�gq9��o��?Y�<�y'�"j]k�C�/��y擝��b�I8"��%�N�Y��^;����fY��lx�U�J�'��o�h��;�N<nq��vx�)�}qp]B0�(̌'z�m�ȦeX�#k��|v'�4�JFq�k~�ւc���bo$�*�ho����Q�*��um򆺺�4rR�O00��;�w,3�4y:���H���.��/�t�����7Ŭ"�Z���nn�����^U[�ȃ�u�O��h�2�#�}���ȁ���q�V'Dl����t��)C�,����n:s��h��L-���9�3�m�[җ�&��VΏ� SAf�Zϣ�Ĵ�͍[~ؕ9iq#ŜC����U�P���~��&�D�g��,V�}6Y��\���V��Lm�
��oj�K[-E�"�����˶	a�q]��5�q;Z��d�xbb�5ΞZ�����oE{�9�������
S���l侇=��wʰ�l����eų����QC���Z�0�	�M�� ����u�a2���U�������Z�BC�] ��U0K��R�у���++-�V���t{�o�կ�.Z�6����O)�s�CY�/y�4�ڧ��%�1�;t����n����-@��s��Z�ǝVn��d@�0߅�3��+��p�a�ފ�������Z=��/;F��8/{�-��3Ntr!�*�Ur&��J��<���~-b��'RS��
�gaO�� iCfVK{��k
�LV���s�����+C�cX�Ͽ�[�0���QІ��Χ�,8u����my��Gg���+�R�.b�"��)��W��Z�4V���2c�����]����Z1�(�}̢x{���>���d	���na=������΍4�	q�Yt���@1>`�gD�Q�w�G@�ĳ��H*�y� D2�O���@e��j��B�|�S��L�RWv;k6E�D�IX�� �\��I��w��GӱR�f�O�jRY������/�\�E(S�փ���5�t���K��}��"��/���q�z��p6�5mܚ��>��?���¨+*��������CK��J{��1f�W<N6�ؼ��=MN�"9۝ײٟ u�J�#�T^�����?��h졑��R�	������4\�fsYQ3ʄ���@�b�i�w��]�3����Q��������V���;�M�D~�t��>,���{
-���9���Y5𜑉���M�&3X8�XGu�\&N��]Bq��$��E���J���-uS�ҩ-�J��	�vS�wt�u_�.&��&��%���}b P\��?�n��=<@���5�+*|
9�m�~�dE4�<���d`_GL�	}F��Z���+��\9����)�@a���Z/7���h���m�;)%��xA������J$��'��Xn?��5�K�@"�ֵ)V�����e��C}ХvM��p]�K����7Y�^����]	rlЇV��Wu��i�s�(�z2���>q�Q~#"��tl �Q�>����!���ԣ�� ���Z5�{�&'��4�62#��=�P̍"���ԟ����X��3Ӫ9�.BG�o��ߪ�i��B|MQUh���4q_�K��'�=���9v��Qj�:OcJ�����ڽ�M�<^T��(,��q*��^#��D/�)�!#���\�#~3{���aL��M�Yx��L���1�e;]��N<5�^������#\�I�k�Uf�ug�F/ O! J�ʯ'�2�ht�����+҂"$sg@�l85�3�&�~�$t�KP��G^e��?] 2�*�#�Ȥ�S��`h�츝�y��l4Z��A�ɱ�IZ�gf����d�����iU#�dE6N����9�ra�d���U�d�@�Թ�|b��_'�w��m[n6�c~1��&�W�d��e�<J��D!���ʆP�0/",�f�dv9�[�hjW�p��K�+��L�;� >��Uk�w�yAͱʈ���Ys����c�:φ��Wo��l��B�yM��W�%m�:�O/����~��&�໌�N�7:P��O{ \��!F�c�@`�-�=w�Q�d��C��������latt�ɾC�%�gk��|�����
/Ph��b��%;������F�9����6����=rF�S��7��LCl3\q	Fg>��A-3ȩF�;ǵ*�犘rǰ2�R/dVl��r��p��H�ܒ���#M�s�4��W�B�+?E}m��Gn������O�6�\k��.e�H�S�/���'�q��Z�ø̶��I�)I�4�IA���鿃�[��KQ����HxU��X�## %P�ZA��k#d�9��:���r��X4Q��-63�B����iZ��5x�/ߎ�l�/R/-����t���hd~Je'��Ϝ�7�G���]�j����4Q�T�����6=��|�%�C��SQgh&��6�KDn놩���eF'�
5k�"u��D:4h��K�mgZ����i=�ҿ���z��n�w�9(.�jL�#�,2"������훭p���3$�"//�s2��Y�sm�����]Dy�k������W�O�����Y����|����{L���j�U>�`���o�+�w�n�y��H@�ɔ8�M���k�H�LOg%qʓ�H�k��^,3~�/}�r��)c�ps��9�e�ؓ0v{�P��u��0Xj޴�~�{MU��K�	j���A]E���hr�#�}i�N5������p��Ά�ԅrq�i�q��2AJ`R�Ֆ�N^O�Ða��r�!A#�	Қ}=͕4=�Ô�ԕ�����@�˻m�0��P��OɅU\�^(A\mWW�W��k�7�²�S���>~�p����ڰR7������GV�_(�m8�V�}>�(NF���)�(����yC�?�	�z�y�7=�@�s�����p����3 %i�j�|�;�T�H�,�D��6*������m��K���0v+�!Z���u��q�� ?�	�C����>(�ץ�5�h���xY�B�����)���h�7?��EA��|�π!"G�^� |������]���	���"����A��Y<����|�p��9a�R6��&v���?n�g��Mc�a��7-ԓ�1Y!�yI������ѭ�x�A����ēغ��2x��? U���I��i�g_��o����I�R���c����e�*\2�9eF�Ng�Yy0hv�57��gp�9�vۚ�G�f=�}���ɑϼ�q��A����4�W@�X���p��)q���FJ���h<�Ti���7�����e��D�w����l�������Qɩ��'بX=L�J2��RO��q���i-#��<u՚(V��`]<��W�"cU?��}y�u{�������y������`��)��Vߠo��&�et��I�Ӂ&���.�����BLN�q}�`9�Ng��u�Ď4ť	|�m�kU�H�6��fOJ�­��n߾[���NOyADO���z�����bg@���b��0%o���h�P��	Ҭ�p�D荖�����"mJ���k�k�O��=��k��b���@����RF�����гݼ	�e����/��_6%�����$S�"+>A����e���n��t��LZ9��1vt�0a�a�::=%�VX��ߊ�B�pnzóy4�`Jq(���`>����5U�U��h�g���,F�Xa�C>��+%�a]8�J��DJ�>�Gw�^�/��~�b�E(��?���)Z�.\V�izӍ�  ��pG��u���s~#��,r���sʮ%���~��|v�O��l~���n�6繝j���ޒ������K����5��Pn���#Ffh�3R�,�����!��(����XN���Z��W���q������0�k�;g��cq�|�xv���M�*���}�ۮ	)?�M	���1}�2����F�KkL�,M1��Դ()���œ�r�,؈�k3�rp��'�S��D_����N[bP�Q,,�%�s�D�œ5̴��PH	�U�q�_F8�L7����(k[��B��~Ä^�7�KR�[uC�_����x�����?a�^O�cpe0�k�ŰiC��+R-ۚ	O)�nɍen+_섕m�	��j�P�w�z �u�B=��A��|��wS�E�ۤum��%֬s� �e���{�K�=5���_�+��7-�sjW�!��T���^��I�lB��{j93��Ip�7�!��s�f�=b����95����f-���ܯ+V���F��J�X�g��-p�y/%0�kH�u�������.)���M�0Z|\~�֟����r�T7�z�*PU���G��󤐨���!S�ˇ؁����י�i��_~ž��x����$�;�$g){zm���ft��#`���Ҳ|���Y��ZUҫ��c����6�b>xIO?��:���r砐�����F��n+��:�̂���+}���qƠ{�G�����ޮ�Y���A96Z=q�=��ӝ�%hˑfB�$�w���	��״(F���d��rs�v����x9I��3��Ȕ3kk��דg^E�B��R)�� q�\�J��߆�G��9�_�]��t���;��]݉��mm�d9�}�YN:���(�H��.$]3��p"Ö#��]<���"aLIF����i#e3>q�'G t���R��d�a�����51K�Z!�z\װZz�9�i�C%'��s�\���`#�1�j΋��J��ՑU�`���D�h+=�d��N�!��ɜ�V%��
B��ώ�˄����΁�Փ"+�g[ʐ}_��^A��[�]Y4�[7jL>�X]Im��^�S5��a�-B�I�09?k���^�R�2�do���+ B�_��Fv�Boro&���o��Q�*O���=D�@E��s���I>}�]���Mh��lXaR*�j$ډ��l&RK���ڢ+GK	ɂ����5����a6��C{��/�`��Zt�s�<���������c�<.o�dR��;o�����n5���4� ϩ��ȝ���mo,s�yO5�,	�'�QE"���Z�,"q�Ԓ�
����g
��D����_�k�ʫ����D?��$����~�|�|�Q�HO�j��+}�P��C�bܸ��f�A�:E� ���:�f��J6��xO�AϮЫF�G��(�m�si6���������ifa6����TY��#�F�Q������ݟ<(�ز����k ��}Fi�͏���1$JF<د� V�Y��s/�G��ad.���sT �^y"]�{��f?��r?U�!��nۼi˱(��z>����xă���WM����,9�a�)��{�� <�:��qKI/����LL�-y��<��3d��~��"�����yo��RQ>��͡V�&�YĄ�s^�I���mapZ�=�g�;��/��f�e�@X���O��eh�	�Rg3�:�ؗdn)J퇒H=����I�g��"{�/x?J����TDL$���־-�r����)9S�(��f�g���a͇�=��ڳK�C���66&a�`L#84�%kN���4Cx��w5WU�M�����l�d�����{�'��!sĥ�}E�ib�`=�\�Y���y�!���x�Z�e��7���"�C�8\��H<�Y�
�l���>��P�}�t|k�N�<�trj��2��������_�X�A�\f���u-y�Ǩ.sG<<����Ѥ�4g4Ւ���7 �pA�j���O����^4�_��޷{�F�Ʀn{-ȲEe�6b��&C���)�p���w�d�g�S;��5�y���e�x
|��� ���E7����.X]��t�r<��ͻ�Q��ޛ�}M)���S���� a�X�V���W$�$d]�!x!ݱ���亐6�%��>��G�X��ů������Yvb�F�1J{��d!d���ĩ������8
� ��[�+l���� ��3����R�E�)IPw��R�ʌ�K��q�wT�}&��~>��N1H�+�B�L_9��L8� ��!d�D���0�jZ/���GW��}ņ%���� �m�����X�֜�]��џb�V��t9��>%T��Y�G��Cz��R�J��Us�eG_��΅z,�u
A�$ƬO�&�y��KrP��t�L�����
wkj�����uv�Tɧ�K'���`�[�yI��U@�4.�#d[��t/��]M3�/�DcN�����]Ő���$KY�1c�T���,�Ɏ{MՆ}�\�@Uc��Ɏ�_���i��F���ݟ��1
e�#������@u{;f��t��͙�8����|)!�h�^-�+�M�&�t6=e����Դ��b�*�*ҽ� ����Y�L��~+\�O�.7J��A��� �-Z'b�o�'�E.fU���R�8�B҃������Ԓ��	B����G�/\+��f�>���+o�T�
��۬s����+��cKض���S��%�Y�L�0s�a���̌l��Z��ֲ�G[ E�!�9�'5�g$��"4��7v�c�"�ƼX%��Q��~_}l ����D����� >n m��;��F�ۅ:f���S%����/S�N��d$s����"��Ի]�iF^����pk ��̬b�6��4�p�q?J�N�+��]K��$4�Ev~긬R�T��UTB2�߳�cFrUփ󩬜}�	� Z�2�u���^F�Y$�!q�0Gu���O���$���v.���B�Y�D� Q��R�FPt	�	þ0�I�b��i�6y����������h����u�]f�fm���l�M����m#��s��R}��^P�������u-y�x�ݑ��Js���tdF�������h�9sG����%��r7=~oH赎h�|.T���{�4�=b�Jr��Єt[S��p@Ջ��<E:� �(Q�\ִ����O.ۅ;*�&<%ܵ�ҏ����+,��Ġ-�����|�t�Y�SԵ�2aY�lK5�FK���Q�vNآ��j8И%w쮋��a�I��t\.���XV12Z�A��-j+eWV��V�=������mp�V��� �>�s�e��QS��J��e�+>�?�:NҸV�p�/��5�K�o�JW�����c~�?�E����R�i�&�Rp� &����2XcJ7�c	n�2���R��@����X�&��eS_=v�Gk8$��
t��j�8!:ə 8$w)�}@F����U�ҁ��J��-�+ODK�ԫ(�~�A���sy-�~�|�ZI���ƀ-�b��&����I
����~(�6�xe����Ov��s����#FR]�%�����UC9@i��}�� �'Fl
�Ԫ���3�m��~��5��ht�I��������=�	�Rs��>�dk���ĕ#�Q�~An����Y�ޚ[�ޚ����qc��&k�3<�k����$��kWv� W��~�*��RM"����R��*f��?{#�s8؜�ޢ��mSk��]�ޜ{��S������#�{Ƽ����	��֠�2�m����ꜲvD���O�����tL���Ѡ���mn(�gKf�n��d|������O(�]�/`+<�Q��F�t�rH��aO0�=�a�͑>95,1(����������$N0�8�4r�1��3l^��"�~�58{GE�¿x�{a5�ǖ�.�W��ru|DL��a�J>���@m�6ڬs1�e��yxZ�
� z�+����$���<1»��Կ��[WQ�����'�F^N�?��Z5Ϊ�(L�)�Bc���N�ɽ��S*�I2���a��@�RLէ�����nH�)2Z�V�!/�����l`�Ӝ'�)Wk%�i*{���H��]�ٜ�VZD�s�]b�d^���p���7�H�IT�)��T!l����8�x�`2�Q:�
��S��UyO�������Y������x���t|B���������,.��A.��d�A�Zf8s�%�VM�[�q�����-xDtX#?����؀�M+��G*ĵ̓_h��shF�Veŀ���O�Rs�4��'�Wi4m�e��`s�>;_7�|B.ڝw��l���I�����W��'�\6���ڹ~%�6��W��w�)x�Ǻ��]	�R��\[̏�R*��H�&�P�8�����O�钱��[ל�*�X��|M�fî[Z�@���D�eO7���K�l-��2�|��;�r�/7D��!�4i�v�sg�<�*�FjEK�F%�1p�^X�}��s�E^g.��'�p�J�'̳E�c5�1{�B������t���΃�4~��(�۹:&#�m^�y{1'�$B�/�uƵ���VE���Nֻ�\Ln��V~݈�b�#;49B�Ԡ������je�3�Ș}v��ð�mo����B�+<�;3e Bc����z�M�K@m����BG1[�Gh�)�5M���8�c��K����ԛΌ�<��n6�P��V�s7�?�4b�~\��K� ��#ȍc�C
�Y1mWe����{�fv��F8f�sO��b�ߤ��T��nf���t$�K�Mf�� ,�K$��v
@�����[9���d|Q��r�s�Ǐ2NT6tBRl#hO[��$l/�ai<"�d�]K�=���:x8x���Ĉ2$�����>��	�?ZhPB���<�=;T�����ɦdK��g�(��Ca�������\L�n�}:kj��dO���?��+�;�[\������/�dT��xb����*�~]|�`d._4B�Qg��%%o��@�	�����~��}��O�
��h�><�csV<���~`�3 r"aR�V�^�e�T�X���W�vB�I�z��M�fW�>N�U� ��|,,XV��%��q�9�,�ࠤ\+°���LCCϚ$p���#��-`�í�O(�u[\V>iu9���j�3�q?-�g˥�z̣'��Rϒ<��>z�'(��`s��
�	��q�	�,�iU�+�֨����C��bm �I��Q� �b��(�!���"�&�	�T��c���h!��j�c�FG��-HcDRQ#,�#lu��$1�zɕ�|��W�Mc�cs���ŽՔ���C����.�A�i�:a�+A���aO���@��?��ͅ�������𕖦���^��C~D5��X�����?\�t��?{���2B�Uh���ܚ�"5�i����U�sO�T�.+�T˷/U*�ڲ��Z�5�7y�&ƍ��I
XO4#GPV��,���z+l�3�^��ɻ��!zf#�t��cq�T"��>U���l\��A�>�8�l90�KsY��
$b޶R�
?�$D[KlN^�}�T�S>����
��f>m�h�Մ>rt *πU̾���y�ML�3�������	��B�J��{4֢.͔�5?�GZ�ྎ�N�5n��}hp`٧���FnZ.ϓJfwnm��'-h")Ξ��
���h��e�i�bMPӾ_��}�+ְ�I��ZB��J�3�n"媧RSk]��k&9��7���+�dP�l��w�����6f�@�[����G��o�s�&_�!f8�
�؈��`x;��Í_�����f�M�q��sm��4����F�{;ȇ+�y���me�������.�Q�s�lS�d�����R΄�8�#�YZ�G�}' 0�mˠ,�q��o��\���-�4�a�]6��t}����^i���0��Eb�~c�ݷ��d�*W;���h�ʐ�yM`�K�-e�i���v���m��x�M�<��k���a�����!�kĩ�!���`�VW�eȐ�d�88WY�و�83�.�R{���x!]z��]W��Z�`���6���������g��Q�w˝��ިmN�!v�� �dĐ���;*�TI���'��e1�2z_Y�b�^�ՙ$:��%��d�=�Ğ��CL�cL�剔�n@�����\��sl��P�>*�'n_���d����3Yֈ'���f��Xi��뉾j8���_{fW�������&���KoX��	ﱡw2 ���r�^����uY�/���%&�Gl�Ʈ�xM��Q�с�$��Pp��v>[��Ϣ�ʕi���*�G���>t�U�|���<(�ɫO���/c���~���|P�Z��ZfD�E��Y�L��+x�3�W@=���!rEdJ���u��B`�i�� ^�����<J�Ӧ����e\�V�%��Ȝ���<�����ڕ�Pр��*���k�GX�>�@��i狯q�Zյ;)��Ä.�dy�lFNO�tjK>&��g������T�r%��C�	�,���<[�I�&��:r�I"��N�3�f �߈�lO�p>�Ӄ��F�ƀ�?��{�F���{h�CLI:�0���C6]��>O�_	�_�07�iCs�K��v����!��\.��d �Zc�Mv�	���g�eut4��Q��{j�B*�4Q��g�"�����RHa��`}�Ш��B&���GcJ
��κ�� y�d+VŮ>�A��{@$O9;2��[ǆ��ע=#����'�男Ѿ]�&�p����U�����$�}6����R�U�ʺ�A�?�"�-5e�����굮���ܹ2��^��ߑ������j�3���|��<5s��e�P}�toY�=��U�X�����`�X�L��m��BX*���h?��\�Gԇ�p� 0��&�:��(f��4�$h<�2�d\�S֭2��O�
Y�q��e�Փ��G8�aP�%~� �G�I��Ϻ�o�XG�v$Ջ�>��y��h�b;G�R@ΎU�"�V۝GJ�q@X�U�Kˮw�=�4��J7;�����VG������}ߖ��c;KQAY�@��4@�-�}�oV��
=��V������F���Y��ydY�e$�?n���9W�{U!��̨�����cтx��v=���q��"첀���8��ti�r�*Ȗ\T�,j!z!w�ѩ{&����d;�u��s��5��][^1�3�n�
:���d�����>R*t! Gp�@ �����/����럯궳�zP&%G6��L� ��N���u�6s���A\�d��� ��\�@"rA�;�N�9��D�Bh>�A���F<�齿.oPPA�H{��M�xu���i�@BQ���X������\�m�Y-MȬ�R�K\N�?��"���QOe����3�ڦ>���H��T�h4�ˣ�&.ZJ���&t��R3����h����0sWDѫ��m@�n�6�?],{�P8CD�&Aa����"�>�����Ш+�ѕZ�̣�D�2jg��m�[%�ٳ�F��b�����m7�Z�	/l8����T��$-�S��D�+�}�����dר1�E�3FE�}e�/�I���P7c��d�� e�z��y��&�y�����������&(��\�5�����i��Q�-���i��c,ٟ�6B�
/.�LQ�̿���\e�	~���f�k�\	6#K�R��zc��Hw	�5-��7�n�:1��^"޳�m7�4
�'��Fb�d���Կ��)>ϟ)ܹ[g�O8}��A�R�G\j���Ѱ�M���?)�vӓ2#�K0o��f�D'���� 9���e�"��3�0��,��e����u�tZ��n����`���Y��c��3�ӣ�X�ەf��yBP��L�x���H���p�M��S����� �bZ��*����c��oֈ�Ys($XO�*u+ޏ�����y�d��4r	�#n��b��Ý���֛لm�O�6_]�xl����^��pBu����8��K��n���}�;��پ��J�C�b�;P*jIՑ'�#�WTf@JbJb��1縩�Z���g~�6ϊw�Nzw�`���4�t��y\W{���+�Y���Us�o�w�O�5�Z��M�+��_�Ӌ�RK�ؔ=��]��X'(fP��	%R$?�-��'�Ո�q+e���F2�Y@W`�0(�D�Z4�,$�����.k�c��9�)��6fؼ'�H���Q��k#�{�0:� |$P~Odg�r���^��������FPy�o�����o�����)��L��Bdܼ�1��D�K�
r k�8���A�W�N��U3�
�j23}�;���0R�#��
��d���	Ͼd�9t�G0� �m�\:�'�)�F��7�3WՑ�-�k�S�<a�mEl�7la=)i��ꎵ��4�yO������-�:B�do<>�cD�C�}9�~��_^ɟG����T��
e��#X����\ucƼ�L�/f�	6��V^����O�/YA'�^���H��p��R��t��D�;I�������S���1jʇdx�K�D�#���K*_�T$�f�BE�c�0�ƈ�J�8�r�Ʌb�O��z�rL,y�Le�ܺ��@y���J�h�z�^"������ƫ�=&�Ǭ���<���h��J�H}��$�XЖc�D��Ms7v��x���3EFpG�߾�F���������n��{)�F+�	_�"����iބ,4�1�к8�rKh5H^jM�z���h� �ۼm9^��ʎ�hO=��yQ�^��Hj[�a�í�������^��n�3=n-��X@���=�2�\0�+�m�� �v�0Y���a(�}D��兊\&�K�T�p�A�@��������r$�󡣳J��>�+k��s�:Rx {�b�]+x�������r�&ʧC��w� ��wt�<��������!��L�g��7��Tͽ��fRNn�i��B*S � �~M�Df[|ߋ�p������+ ,BgM4�<$�3�3�%͔��&�ʨ�L��&�<	��qț�`rjP��5�n��|+��u(��Qg�Z5�~�-���\U�7W8��L#�m�#1�Rq�L�dOu�Ϸ���{��2~\�شchVD8#�@���Y0G�P�SR���=Uy�y,�"�����%�������� ˚�k�:�Q�Nۚ��`��9� �}�KU�N�p��O^A �7�4�nZ]̐ /%x��+�x���g��H�8����.�0�f�{O�6�P��b��͵�[<#�����pCu=�ؔ5�HW�o�+:�L��m�l�;L���)�<?
�%j=X	k�r�P|��JNS��|C!1D2tz�����: UM~I �cJ���VSJi��?�w�)K`�fj��|�FP+s�ww+�����9�x�B�/��9����w:���K ;�����unal�~p"o�eH>�HR��G�������o��AQTlxZh�jm{YRn#��s,yb��8<�¨��t@W�U!��I\G�/��DA��(�״��ђz:]�Dx��HSh�0�F*�,�e`a&oÀg���Eg_��@�r�Ɯ��c��A?챗�e�WJG&hf*{��Iêj���O�&�]*��ױ�ׯ�� b�����e��;=i�ۻ��F�嘍O1�+Fqqc�#�qJe�EH��X��M!Adͼ�S�6Q�t�i�o���Un�|���S���ê�ٲ�:���&n?�Ū�.R��k̲�+�$JE�G�#��xf���nE����REW���sB��
�M?���]���te�ZT׍��Ǉ8�.�+��}��k���/���k�B��ش҄���U2L�?|�> G!�rn�I-��w�π�D������3�fG.L����t�3�U���R�k*�g��.����'�!Bq4i�&N����;�QD<��1�ޯn�6Q�o>L���s�&�m���fs�Uln�aV|w�Aב8r�2��	GC�q�Dh�>O"?����r�TW�=���E5$��>���y��Uy�Z�C�ؑ��8�{��.��{r����Y����9LH`�]A1���4۬i�x�㝐�!��_��x���bm�_5h7��c�#b,"!3����R������t��h�?Fj`LEe"�c��x���"��#H���xm�7t`;�݀w�K\�ت�ϵ��� ��͈Ff5,0�)Q�ȣ���N}�<�:�����0�z�Ŗ�/��~xE��3�?��wzJs���I��$���I3z�7��M.�^=��;'Տ�hУ�kِ���TRcJE��\��0%�Ȑ-r�g^I3��'1a[Q�ƜW$�jlEcy<IWFçi�}�~	���֒���C��lCI@(�ꭝ���[���N��s�p �L�j��_^ă�P�I�Lk�����}�j��E�M�¦��;����T&������l�9��Q���ݻU�d�Gmd�'H*2�h�fT��`�[�}�	�ӣM=c�Z��B�<�.��܏�ͦ"�8F���聎�Nh�J���[���7�*O~-�l�6uۥ�A?4�Sk���&�ڠ�3�kU�U��a�{��
�@��L��z��ψ���G���q(?n�+nEx�Jr�Wn��;A�o��[����u�P!�.�V
�r�m}��i�N-���m�?� `��F�D�3��]��j{o�PU��x���l��,�@�����/�>Ā;,5|a�ض�H>���VG@8���,TH�g-@���\|L�5o�<������n�m`ɹ轡_]�&%>��<3��<���¢��m���/�(�S�x�|kv>O:�E1b=�{��%�]u�0����Sv:�Y
f>�)8�?)d\֭K�X{�Q�Ny1ܫ ��F�?�y�͈��|�:2^Y�^��ŭ�N������zk�Ԇ��{`0��0:1oV8x��^u��Ǜ���%�e�����ƈ�+F~|�~%�8���Yne�XNUӻW�0�����}L,�����0�o2��V���.3�-(u�O�J~�?v@�)��>��ƹJ�������8��Zg�W1;�P��Nثl�(fc~�Y��3I�D82u�oe���߁�����䅴��F0,�⼹��#�]��5�^q�7$8�c:�����Q,V��5��AL��vU��2����y]Qڌ��M��(�Y�'Bs39ˉ�VT��
�;Nv�3e����"ya��R����d{�+�����`��w6@111�jG������ݐ.���$�7��*7��4��L�����5�c�՛�~5Sύ�K�Z��Ǒz �Ι4�\I��l���壘5y�X��D�^�M��a9Z�_���X]�(��N�lx�=�O�w$���$��_uL���W�6Y�ܩ�v��/���w/s{B�7�+�������ȴ>��.���������Ƈ�4��f?���4�+K\kz�=�^Ot�i���77B����t���M۪NJs�3:�����aԅsZ"5Jc��J
��˘Ր2�\��m�7�i��$�XoǢ����0�vP�{�\�`5(|6 �?[����ҭ�^�#}x���=bV���F��=#�v��a��)�G'ź���0�ڹ
�ߒ���YB���U��g��_B6�У�$Sb��zYPJ��E�q�Տ�B��0eq��V'ψ�6g6ѐP=�[}mya�|:�a�y@�Q1�O>�F�`73��ҖY�Ev���RZ�C����C!�� ���{_%
Kp�vc��s�tT��r6>"�g��(���-2�}���uO�HݭWu�̒���KOӭ��} &�}q�PWy����j+�,�jh=����|Ҋ�A[Q�"�')m�9�qW����Dr�R�v�.�E=��7�ZX�&ʵ�(�9�k�Cg�%Hۇ�xԈ3��T�IX_]�8�G�I&�ȿ�Qw��#.�-���5kF��<��#���o�;����,���S��
6�S�6��d�h��Ui�d�8n�+8�~ARe�<�X����`=�j#٧=�w�����\��8	DBe�x`b�E�����iY�"}�6�a1u�s�NSq�J�ıSlUC 酕�!��缎�	�g�:�"F�Zk���X�M&L5�1ˈf\N������ܘ�K�tЖ�����cĪ�a�\JK���!lжa��C{�-�cK=��y?	e%�����i� ���K���<�K�7�VA�>��&�ˊ�A"@YH�zw�<;�=�ag�~���4%a]�|�5����4�r��q��hֹ�'�88 O�.��8(��V��4YtO�	�k&���K$t�BxO�n����*�s+A�x��N!�g�R���U��ʒÒȥY��;������K��婺��_)������S��24��vy�=���wЮF=W����V����z������Ѧ�^���pa�T�L�ua�/�D�|c6�:m���<I؀;y���M�tܲ�͚�5�l��w�
��\0.��{>8Qą�C5sw��x��U[j���n�?�X՛�1�f�N;�yHMtG�D�c�]A��f�a�}�Ⱥ1j��ڌ�yu ������*M9�v�2����Ssۧ?n�=LԔ� IA����5}�>ٝ~���� ��"��p?�~)Xi'<�-x���<2=�:���|�G�z��E��,�q��^�j����a���_�;�vB�>Sx��?��
����e��Q&|ӳ��o��2��L��ӯ�<�e)�Ǻw����7�$t���ߍ��`#�\M,�W(�c�f8��������� (�W���o�(�e�&JWc���I3�̤�@8�/�/Ɲ�-�Bhh��6�::E��<o�H�!B�@�&tN�u�/�`H/K���yŮ	w��8tg 5����:��|��gр�~�4��T�Yǲ�C�rي�2�_]Dӕ�{��f=�y�����s�q*�Ӿ�`��2�PwTv�y�Fl�+B0������f�K;`�+����4Mia�O�g-��Y�LQp�E8-�Y�{��u{<�5m$�8]��%�2J�[���#��V��by���ݞ��pX��4^#]�j�h&�a
�i
ώ�Tx�U�YgT6���!'�d�D��6���T:���� �F�����A���8&^0�܅V����u�x��?�g:7T�e�Xu�#��8Ě>���B�~��s��v���t��X������]�ĂD�Uy�Jnq�I�O�pi�;Jt����%4�2PPL�k|W/�	j�F`\��������i{X��X�1_�YͶ8)W��A8�\����
j�n?[�9z��ǂ����6����qPZ{Z�K*Y��ȵ�}�,L!]*��=3����K|�6oH�jcq�!2�<���	Ů�˲�u0�ӿ���c�������g��W�|���݁Ɩ�	.��#��/�Kd�
��fz�>��,���/��E��/����G�O�bS	(�y��c��G�����x�(M�	*� �@��^F鏽�#u&s'��?#S�#�'/�� 
\`M�FFG����|_�+�^]n�tJ���-�
�p�ؤ�K� jX*�����>ܾO��6�,�Q���+{�r����Q��N��Y	��i���;���%�H�&<H��a��H�,���>�%�:��*�à��h/e�+#�
,v�Q�m}�B�i5R���Ώ`�)�_����V��ڏ[�ʹ� j�͖����sA�lF��x��JN���5`���5�P�l�'�R�e΁��_�亣�b�.j��z���F����>U��|��D��\Ƥ@q/��$�
�O0�1�ﲽ����r���
�/
�Ŗ�P^�3�z����?���m(HǛ;9�Ru�.��#¦tdSZ=E;�|��-L�d��}��	�+�W@$U+4�S�O#U@LVV;�z�e�$~h`���0I�,����n������%C�N�kz�Ar�5�<���X�]�!��HZ3���Q
�C�%��)��<y˝���ۮdu���������y)��Z>�?.����m�~�)��ϧz7"p�+�:ϯ�m�x��e(�z�hxt(z)Fn���B��2R`��O��	n��M���r����-�����,*�0>M¾֯��d@y�3�k����pS�-RO�b���{�İKt���S�Q���g1��� ��4�̛P�M���Pv� �.���ѯ��r�L>P_�W��	�xy��z��$߬t�h���z�����( m�� ������Y�y�ԏ4ww�	H_�S��[�5�"�vA���z�	�X^���\��z�v�~�6]�~���mh��>�)�e��D65���v��60�p,@��uzNʝ���A:qQ�pg�RV\�5h1�pt��a��~�:ڐe�礲� ���U(R.c� �x�&W8\?P�K���I|1�3[�Vmg?��i������8����rh��/����.��i3��_����s�o�6���:f���<Ъ��ٽ&�!��ϫ����qg�P��vY�94VaRi@�F����3_a��r��k�NŔN0����m�w*���6	��+��$`Ai��Ҵ�,��#����¿A�n H��A#Y��8
��>tsK��t!��{y��(�[��$��m[%Ǯ������.���d����wHQ��[;+��ܮ��
ØG�����Ht��V��K͜�O�TQ�R�n�J�	��(P�?]h�ܬ��d"�_� ;�5�� �*j�p�Z�
n��Aٲ��H�/���vXp��h0�v|��ɥ*ċ���5=m�7x��Ȼ(-xsc�g&�o�JU_�_
��e��@��*j�����/u|>�M�^�%�=,D,Z���PB�M�KGۂiu�<��Hr�mюY��-e^v�Wł��Y��c������c��s�h��U��4�s;��H�IT�<M�|��6�0~��§���2�#�涶[Ts�G�O�1�ŰVNL��.��(��ӌ����b6����B��Rg���I	�"�b8n�eΔM����p�n��z�l[�p R�lqh�l&��o�8`TTe�`�]	oP�)C�V��CSA^?��1���8[^���QA�����9u]����W<�k��n9t����'I����_�>PIf@�~��y��e�d�F�O�kS��ܨ�i���)P�d�
�=j�� �}��͆M�E��C~4lm�OC5*����T�'$�6�!1U�v@]$
:�r�A>���W�oBh��k�'�P�z�
�H���Λ]&>��Csp>�C����S3y������j�Cr����X	ro�t�!hq��"���
ƴ6��#�g��x?oJ�t��7UT=ieQ|o�*E��/��	����Q"�H�V��U���U2J�~]!嬢��S���:�N�����r��o9� �Qj���~�X�_�y���E���zb�����5�5g��L��#r8����mP�*wJ���.J�{P�f�N��������@���8�8c5�8�
�ee�{ԧР���V9�����&�&�mC��pA�TG�M��9ԍ~mt�+/7��>�E�@�Md��J���iE�(GS���������p��r�Ł [�F���J��d��懌R����WJ��+ܝ��x��M����	L�n�~��H�P�ߠ�����~��=�Ƹ"��h����P�<�ֹ��[�4��ёLwY�Er�ۣ�/�j�q~��x.�����&U�a�w �Z�#%~���� ��f��ԭH�'չr�<3ÀC.D,�$�ށ����$(�	Fz>֠�0|��:Y�K�K=ڠy�M�|41�ձZ��W�]�<`<]�!A��Ed>4���8���O�����(@Xߏ['pVCe�����|���:����":�}H6VH=<_����n���x��L����n睅`\t̔ie[�����4\�ö�m�Wl�t� =-��s	%�;��~(����1Ɏ�&�->j#�XVʺҠ������=g~�͆X�_�����Yk!�W�&K˰r�C$>{w����:����N��S4"��<�Aq�Q����g�J��Ǧ�ޫ2u��p�5��P�L��=c3��8�AW��4� ٩>}x��k�~�f\;��cH�ȳ� �=w��?�Y>��a��
�ec���{c^TB���n+>���+��P���	�j�.�M ��@ߕ���pH�5$l������*E��eg\�rCA;�M�Tmx�;A �ɀʇ���Y��K�x�k��D�z�l��>�`����'=P_S�2vg�u%6�<�+�����!�ic���pF�%�v�q2��8 ��lm���z�&L/�(f�u�[s�ǋDL-G��AUY���7	�w�H>�u0����+�I,-#E��蛣��"�\m^���[.��b~�O�J��l�ږ�z�i`��K, ��ʠn�ۃ������6ua����8ww�S����H"�>�+��4��|�q�³�~Q��!%^�Ɯ��vh=�_W��4=&��ks
<�RH��2)D��j_Hj^�l9�S0��ո�)�t!D��n�M�&A��S�T�� �zũ{�n!8����gO�V�r�$�5��v�������x�R�Y�ˀk�9�0��'0���q�Q�S̲e�[���x�S��D��f�/f/ ͱ#׍yD�e�ʊ���u \�ѹ:=���Z���J�D�����*2ev��_�}9SL^5������@�x_Zޡix�Sf78YDȔ�f��	j{+L�/Lpc[n���[cIx��mb ������w�D����|�en!�WJ�_bBܱ�jh��l�����s%�:�K��e?�Bn�������Z���w���;�j��֨�l���ٓؤH.@�tI��R�=�����ː��h����Ḡp���ǸS�^���4̀CvE�6�_�t�ۓ;�SNt���g���䠕Q�H�)�}b{I�J���ƌO�v��jX��e�w��v�^�s�F��~����r����T���H�1+�����Os��d�y�x�52�ċ����pN��sF�o[���zwQP����~�f�U:Q��we��
�}����d��(X�[�����tM��L���YUU����2�.����I�Ee\����h
X��6�W �Cl3��Lr�,�#��t����M��:�όgqW�*LʋJ��t��V��J�6so��mѡ�N���2r��Z@ٶz=c}��,��re��$���8��'� ��`b }U���D ��w �P�`�ohpns�������ɩ�]'
���*�.�)D=<�Ooo-�4~��H��|�x��!^�n�w=o�:	DÁk��oG�P^��@��ŝ���o���@=i�6c� '�0�%���#W��ka�y���]�ͅH�:o+?(
}$;���L7�k�}>#:.e��w��k��zh ¡Z4w�D6j���a^���cP��F�*[<�����ޖm�7�$G
� p�gJp��&�����\|���ȭ���<q�E��()P�c�]U���� ���;�����L��mv�WoAd(���ft`��Xf�S�G��1D6oɵ�dJ�o�'�&9�j!,���>��� �n��k�Վ0�Z�^�}�,�����	�(aә�QƄ�pzXd�U쟎��y��(�X&��r۷T��M7�ıA���C�s!�����h�C���L����A�:��yO���`��-�oW<�8��\�re�S<+k�u��9ev�^�hM�"]ܺ����M�_�R^A..ݼ|�,g+�p��BĔz>�����8�2S��:��ѧ����~�Iy~^N"��+��>��+������ĭQ�_�T�%���2@ p�c2ıV��%\��,����o� �L��Q¯��UP�6�˸"OY�)���<:�Qb�'R����30ݏ����L%�����F��%��(�
nZ�������>����.X6Z������x�֋��^ ߎ�A��c��ӫ{ɹ�K8v�)I�m0�{c�G��O��it�d;����s�����j�Py����Q�Xuh���	��Э�2l*Gzz�2�aYUC����12y]��2Α�8l�:��o�Y "G6��$0�a��t�_v��7ΏUv��4i��U�isYs����wNY����r��`�
G�.���
�5e�FT�E��_b�-9,'��W=�|v��08ඹi<łx�.6k���#���`���@0��x�B���aR;g��Ue�|-<*Ya�Kc�L�ɪU"n��.M�h���8�ce����VfrV�M�F���]�e��,l*�G]��騮��%_���s��C�y�(��"��o���59�o��A3�/��w�� �7�
i�M��Oo,�Cn�o�wvҋе@��5�F�ƾ{٩:�(��.�B�D�X��DL�l9���!��� u �a���	yS����%�����ΧS�5�il��@a��/T�U�vj���i⣜y%�����&�3�
�i}�~3���m]��E�9��쓬i��b�O'D��S�Ki^��Oms�h���?���u��j�r���.GF΋�K̲c����~��g���ʩk�wgvH���S~A�5z�cuc�㕑������%���67��@Q[ֹ?�G(b�鵻�=*��ɯ���:-��G�f��&�u�Q�V���(j"���$��T�}�� B���6����Y+��������^X���k���b�cȖ7��0vLP��i�#Y,Ww#�֎�̓ڪs-cq����'�$���J ��E����y��[���:Aa}��Y��۲#%�c�o41�|,k�g}I��Γ�A�`�L���.:��	�zw1�mQ�
�k�h�{�1�b�0z\��x1J+����E�y*�'��d����mBL��]Z!On�Χ�x;��ÛQ�Ŋ�q���6w6կ����pϒ$%��xj2d�t6,�wx�\Ԯa�)�Ą&���c��#�^�f�yT��E����R�>�B�,��2?݀���.O�VKH� ?x-J��8ִYm:�ʩ$Z�6[���v����Fb��p�ﴺ�:��()&�'��)w�ZXj�BB��r���5�.88wU��=�J��O�>��h��3�{*DZ�������0
��Ѫ��1��*�M�Wm�@ !�8@��r�g�]�zm���������Ӵ�ȉ�sB�",[��_0R(ǿ��9�Cn��2��� q�(�J��<{�W�4�gy��sK8%;�����Y�I��'���uW�����j�j���s�%�Xg?Qq��1Yh��)�Ҟ�2_���p��Ķ�`��N������1���ܠ�ey�-͊]�3.Ҳs_uZ���>�n�?����N���|��K$O/�I޶.2����w���2�0�����i	�߹V���i0�
������]|�����/����t�\U"��|�����M��;��Q���n���&��Z�o�oE^S[t�	�7���Y�Хk�d��
G�72x�T�ۚy ���>��$��L�N�W���BE�k���iJ�37D�� u|���.���I>/ز���w*a�"�I,6����J�鼩Q�}��m���^��6m��?��D�fJ;IM�yE�s�utna#޸�ym�Dt�	�
��{�G�.̦��p<�Qu����wO���K��]���)
�3�Q�g��9>�����Z���� �:޷4�BPp%,YȨRz�Z����K"���]�<��0�B/��w�sT�d��6�o9�u���;6s��xebJ!|_��B����b�	ϋބǢh��;Ϸ�<��P��D�$6V��<<Z� �*R���Y�ÿ��lL",ۗJ���5����c����QtU~������m�Nx�Lh�K���r�D�4�Bw��bqV��لI��?�OD���f�̉>��a��5���®��ƴ��������Cb~1�#��M��)39�'���t,����QE?���ە�@G8�U�ˤ�<2�G�)�3JK9b�`ѕ~��#�F!L�s⊻�&lz����/��	a)nk/��s l���v����}��G��nu6ҍ�* �@��*�+���G�aj����"Gg�bt/(]6��b��t^ʸ�a�Ӝ5�y�L�����
�l�j�a[>�T�Ļ}��YjVIg#P� ���N:ӳ��D�{.�(G 8t�[�"x��%�L)�W�M�/˙��^7Eye���p�Q<�^�� 	3]w��n�Gk���җ�����3��!�C�����|6V�^�-�}eB��݈�L1�:1�`�,�E6H���3`m<K�[g��;�u�Z2R�+�[�fh����j��ia������Ψ0@�1�e�E5z�?f�qS�,I��`,ǻ�P����y���S�K�^ ����H����1�D&�ai�;c�C}�����X�s��h�XXf�(9�ñk�r�`i�]u
�\\"�n%'2�O��yC�',Y$O.$I��1�g���P��>/�5�E���U`�9�Юtz5U;��|��-B�hi�ޟ!4@fq��ʒ�&�3JfԬ���3�J�$��� �c��-�>7�9�	!ů��{����矀�.��T����ۛR��b�6���˴F`�Vi�'��	 iA�(7�[W"�w����Ǿ>��?�_�ԡ.�.���X�U#�X� �c��L�y���;pգ&O�v�E���x�3'	Si�3��=%����'v�`ZF�ۯ�e���"��&YJ�&��E�R-�2���Z���Z�D��ܘ#�0�%�*Ph����Y�-S�}r;�^e'i�#�N�Q��c:4];K�Leg���5J�O�)�������*О[���%��Ԑ"|��O��L��},x�s�b��m�z�%23�Gю��ev^>��r �3�$��n�*�T�@Wmɱ�!f�/�f���D�X�$���X��5�y��������`��T���i������n˄ҧJ(�+�5^��/�K�'�:t�2ֆ�[6���a��3N0MH�7jC�3k��v�_���{!������h�n=ǻ��՞R������sA�Rr��Εr8qȼ8��}�zبTv�6L�1ۯV�ܻ�O�"jE������M%:!�63W�"�P��w�g�
do���m�\���i��65�D�̑�q��[�Ž˦���;������EZ*�j=����Ib0����WG�����%��b��]�P_���}_[L�����Ha�U��"�]Z�v�L�w�C�|qs�o�2�.��A�C�i�it�TO����2@�X�Ɂڕ?r��ԔW/8b�����KI�;����{~�D<��_��~�+�mP �c	c�E�㔖����]o<0�A����i<�Y9����.3<6�l������A�%�i3bwK}��0)^����.0�����o vط����Gl���;t:�`ާR-�]���t]u#܊�f��s+�����3�D��:��P�7[_��w�ʶѩ�gx�L{������L�U�us�Ư�2���/�W�g�Y_�w�o�f2[��F��������\ٌ>h����0 ��!���?s:��vmt҂(�8�.��N15Ç"xX0���*�b$"�6����.��6�ʫk&�!h\����}kO���=s�}ƌLK�:�M�n�Ԍl�ȌM:"�d�������=���Ʀy�m�^�_�5���:St��v�Y����[�3I8���PBޝѸ��h������z5���]5�L��^��e{i/�`��UP�C�� ��O]�=oi"�����f�ɻX:�@�q�+`R��KMU�S��T�,`�1� w(�����*�UO�N���1}�P\���ձt���X����?�b������� ��9�GmҦE�w���oa6��/��O�j �'Z@Y*�7���C�*��P�Dܸ��j���b�aHq���JqĔ�.�K"ܩ�G��(ы��#~�Z����8.߇�gȽ<�]Ӌ�� в����D����AN�H��}�))���}}�����N`��fl��I�/H6�����%j)�ʟY���T��PL�R��\`O#�n���o�34�7kV�y�wZ� T>&���LcᏜ��#Fޯٕ��48�1��bqI�Pw�n��������h��{�i���+.a��x�H����3��fL�Iԅҏ���� ���5a3�ޘ.[:+��w[��� .֬���\��	ߩxRjn��i�-�~y�Ah���Q,��gHeB�Gy��5/*�"�l?�dR�襃���֩�6r��ў<�}e睲��_ �-�յ��U�f��x�ﳒt�i���y�S�k�D�ڌ�PF�yLP1-cr�l����7Z�`'�G��u�ߞ�w.�t���7Y(twT������+~���'�N*�'7��N��g[c@O��v��,��e��YŔ�uI�KEŃm�2*Z�5�����4��I.P�`lW�S��.��x0�=�N��KO�K�(�3��Z�Y� `$�*�KB��A�aos^��lJM9S0Sc��������o].���0"69{���_v�k��Sy�I����x�]K��t��g��!{Ζ����t�K'NΈF��y����z$�N�������ĩ�&^Bm8i@\vaEo�IS�ˇ�1���҅uz�J��,�f�_��&�w�ݗ,.ߴ�O��D��<&,�B����gu�HV7�E�(a/��3=z�Y��d�>?�Y�@��g�U��u��RQX���c������r�U������0��X�/�S�bn��?����fZO��a� �?�q��ݟ�joK��to���_R@a߇!��y��'��0�{x�{���D"'s���3�I�3gӹƃ����(T���[Hk��mhR��(��ĉ?^�%#��j�(��J�9�V�2�r�ٜhZBs��F�LԬT��g.�Oњ��$��Q��UyD�u��%形y�NnZN8�ڙЦǴ������H;!��꫸mԅ����\E	�@�6��f�4�5��W��s�)��G�5��i9���m
��{4�z��|)���*7rAE�<Ю��z�*4�g��e�G!���mZDq���'c�覷�	V)��=�՛�]^:y�Z8�'G�M]�&��d�� c�i�A��lϔ�D�s��'�u�[���r޽�(�ca�j:_֖R���L6�?��ޱ��[���*��t-Y�V�?>�\ݼ��E���.7���un{|d�4R�W+��ƝyK��+Շ�S!�na������6~�o-̟"I�h0�w��x�R���������t� |mL�T7%�u���"�
"��<_�e�s����@x|��2���ҏ=�sq	O�CB����1��[�E"��?~����ۯ���6�+Mk��kW�NTeQ���O�w�q~�g�뒕�:m�6:cD@��?ʘ D�R�I�j��@������ɶo&���V!Xe�t�(d�ނ��^�RT���Rt��=�p�BR�|}Ŵ����D�;q�g�5�����ǉ��\�ٸ�����V�M�,�H;9׃���tj�߀�
S�Q�kp�.�<Qd~�A^�!ފ~BoK���#� :��.O��ja�(M���m�f�`}q�@0D��TWw����#��p�|Y�D�p:����0s�61��s7 b��K}`���vJ���b��_�pA(�p,�nu�Q���>�b�,J���@Q+�yk�T�<�����+:�lEv��d�9��Q�o澗��ڡ(�Z.ǚ�7�'�Z�8����]�BՌ$jJ�v�4nji �5�ǭ�5�%F��r��>G4�����NY
�&��)ܰL�A�"�խ~���\z#�3 �������E�\��^2����9v�l�5w��u�<RZ$�������k���o�MZ����u��P�E�z��>5)J�� y�$���7�q߰�\u�&���Q��s\�A��G����C�I7 �c�k��M���<��%�닶����)��R�tuhm}�-|�cCKc�S1� ੾��S��A��V�)��}�y�Ģ+t���c��v�YG�l}LO�:�ϲs��M�s��Ǖ��hLмg��D������E�����^�9�Ø��.�ı5�p:�kPU���V�\�!���AR��Q��OBRj���{��R�����+8�ж@��tbh���~�jF�puCLӻfr�߅h:O�>��xs�ՠv�[l!�aq�;��wb��f�0����d�`i\�c/H����%C˗(@�����8@t:��J�Ur1�����ua86K�XF�]N&��w2Ԟ)�?*l�\�BX{��k�cp61�t���cƑ�A���F�A�&��,]�5`���H���i�e��DC$D!	�M��� @�9��"���}8:�.W��B`��Q���/�c#>�j0xH��<jpͲsG�u�f_&�Ox��ݳ�{Ez���O�^{W?鲥�&��ؔz��Ԋ��mE�+�aQ�ff���Bϟ�mu��J���#cS��^\�]��⳴�7��x�ví��6}���8�W�g�-���S܁w|��^�S(e2�9Y*~&�X}܄�:�^:y�s=o��i�ƫ��[�X����E�qEC.*� �-� �m�w��{�}P���`W��]e{I�9?#�=���
���V��hh�ٱ�us�x�u.8)�ped>霍�2|�U��-�Ҥ\�j�g%���f��p6kL]��ܨ�BK��H�2�yg5�
y���
R���� �-�H~4A;�]�F1\XwkV�z�Y���oƲTa�C����\����3r��
��Ǹ�����h1�ԗ��Ȍg�[KM����f��b��y�K���,$_gF��^� %����VP�oqӀ�1R�+�H.�)�rW��6w?<�4R[f��n�r�Z=~Zd�і2�IK���6�YG����	���ˁi(��ۏ!�&�1!w��������0�;|+I�v]�]l�Ц̷�{��4Od
MRպ��dQ�/�Ӏ_�c	`Q���oݱ]	��HXH0*��z'��x�D.��ٴ	��ղ��|��/4�YR�_������	��.�؋�*����T� }�/�O�9Mޯ�Jp�����)<��_#�z���L^t��*i<b+�O�Ui׮�F���4Ap�d�g���S�vRLT2��h�̆��.FV�B�֋�ɜxM�x���_L�MD�(�V#h���g=A�v�,3[�%����QGlͩG�v:��|~�>w������dAI���C���P�V���U��'O��f7�&��,�cц.�&.5�l���33n�[}]��$ Z�ezS���4��E��9����oI븴+�X��Ĝe*���3j�gS��?�@!�OYD]���ڥF	s�O��ka�����>x/�(*�K/����mIt�Qq5qj��wh}�<g"�ӎ6�|"�5XC���q�&0�O\_�>hŝ|�J�Y&�����.��s?���B��2%�E�_�=����v���Ka0L�S�J5EI�Q�{t�m�^��n!]���;�����P������z0�m��<��B)r��	������7D�` &�!sf/���U�r�o~ѿl�νU
�A)�%j񤥮��#n
R�[đ�ebȍ�\`޷���l�=���:�1�R?�i*S� �^UoPi���9T�{^#�*���?N������w5e��,����>���j1�憪��ՃD�L��Z�
e	���}�n����J�fd �Z7t�*[�9x*
�I��z_#(��?�@����� ���N!���@��v4��8g�dU��WB&n��wօz�r�\�c��D���;[��5��\6��|��h�K�Id�TT-�}5���;8NMkȹ���(ܢ�WU���2��-�'��Jbf���#��ݜ5���70`�c[����"��>����/ت��z�y�+U��ưK�\��pL��o���G���P+.B�Au��]Nc)�]���s���p�9�V�݃;�"q���_gK0�����m���p����Pu�l�z]K�UC�No��;��e�Ѓ�>�rk@�O������㙙��o�,򊿜���S;�5�>} Z���u���Blg���N21ƍ�� 9���D��G.�h2ՍTm'������gH����:zߟP:��������N4��p�- �	ǸAe�@\z� ��Wma+��G��Z@|��.o<f�����>vi�`�l ^����k%����q�O��Ii�pi'M~�읫� �����s�y֘?E_9�ɪ�#���/��;�Ӿ��W�!�j=�BD�	Ѝ�
�m��--��3���?�ȺXS�NQ�T#h1X��0G��cv[�ͣ��t3�O%Oi7d��W���IJ�Z��q�`{.��������&�ϭA���������F�ݥ����BP��)����Tܓ8��$TNݲ��0Pw�o4�!���ޜ%�5��a���z�������� �H
n��	1�hMKDJ�oW�Y�J�z���AHȘ�kW$d����XG���ڲ�䶹*6>��� �y��yz]΀���������k����=�#�^=��3^z�:>�_gWks�r%{
R\�Σ�C�f��|)�Q/&���Ǧ���^��o[������
�U�5���,�{/���%���5����y�w��i	�P_v���PdZ�
�7�$8.�!`^~�q�������<��i�����3��3��JjsЭ�;IۂNN>�״,�L��W	�e�#�[��x�/6=ydr��|>�x�#�%b���B�:���M��E�`"c�3I�c�Y�v~�����q�X�����^}���ic�ʐ��V������h�f܎%q2�ZG�3V�z�΄3`�?ƹ�kG_U��p�EG���tb�cD�k��F܉�qRe�*��4������e�%�8iAs�����q�Z�eK��eA��~�Ԕ:�\s���e��{�f��n��B�J|Q�T�W���[��iث��(�|�Ʈx��ހ���G*q�`2���`_�o�Oں�$y��V�r�a���a q����l�K��=w�7��7v�)N�su
��-�"��GhG��')yfpɶ!�=�'@�D��C1
U�J�eM.-NC?�G�]B�%�:B���&_U��,�J��	�9�W��"��k:�j��Y�wl	ݽc6|��Rg=Յ��uW�q���1@d��L�?�/�K�M��ϼ�"�RX�i,��j!�42-��ڑKU*�S�x�a)�n�w�҄@�x�7x�
D��E�y*#Iq����՝Z�����.���̿�j�`�X��޺���T�[<	]~M���QrE�6�`���,�5Rn���[�
�Cc�������k�[z�Z$�jY�.�*pZ�!Ϊ<@�x�}V�u�Fp��H��B.���?K��$�0hY"��k�P���v3aӸ��h	 0�����2׋(}��oR"�%�6{ݖ��M=ݛ��C���	BI�+�C�G�5i��/�%��'�M�0TU#�;���G����{ �����ª�0#�D�{pz2���G�t���a�rF�4��b�<���LH��}Q5BOj�VV $?�mo�q<`�� k:S��Y�;�k��c +8�A<g�9��퇚n'h-�G�����Љ��"{ޙNue������]�?�0|���8H�j��_ZO���@���ߌ��;#��)	�oҺ+V�C;z�����\G?�\]�L���`Ғ��dc���.�Bq���Ȟm�ǩ�We�����`:0#RH�?@�*�%q�y�4�"M~�4� |7�.l�|&�yɱ��P�ݯ׷>�mQ|7�V��4BC[ˢ=Ey\��]�Gy�縑��2�Z�2����
}�qISu��e<��M~G�m��7H̏�w��������C�:����o��P#��K��tUQ(��β_ܩ�&7N)$b�؝Q�ʙ2�����hKx\�I�R����)��rJ��#k�U�4��6�`Z��6vV�0c/'#���Iqr�����[ ���e��k A��>���4;kE�R;��6�9n���
���;�?ɣs�E��DR�����]g��ս�b^<����}/�E\?��u��'���e��*ȏ�͘�=4���5(P���`@9����j7���;�[�=`��k�x�m�eZ�O�$���L��p�:*����_hZ1㔨���#��i���YQ�J_�¼�B7=�9��bw����e�?��B�|�.m�J��[��1��&a%4p^E֘H��<tBɗ9P�3�b��ل���r��u"��6�r���*��<���_NIi+6��y'����]�!>�; �wXO_3d��9c2Y�/�5ǐ�s#`���G��,�K�4$�ۇkV֮E������͓���[�mf|����l��L��k�jCn6��5uu`�R�� �\txܩLw����_(�"���XӶ�J����p�'Ol�K�{P\�8ї�I���/�G�Zi���B��ܚ";���*b�9P���O)��=��p�[��W�N��}��&������u����~�WNy���1��Oz��A5Yپ�L�� f�!�r11M���j��P��gl�Q�r���+@�n���"����ou�mWZ]�����^w���9�2����6Fȸ=�P���[
Oo��M�ѣ�݀�WZL&?�@ ¼N���Mf'����y�
���,��p����	��ȹ��6�����E���d{�\_%���7S�k�7��M�&���St���ֵZ��޹������6B�AذJ��1E\��U��g� w~ݗB�#�.�3E3�� E�����)�vn���n؅誽/"T^!�������ip����j�@}�p��O�f�����Rbr9PF���w=K���A�8[��C'eE���-*FYGsǰ�ڠ���RE��j��+9�Qu(N�jH��j�w�~E<�l�4"�I[���@l�ښ}vlTBø�p��]����L���9��˯�*�:��kf%�����q����}�Ƶ�>^��B��?�飖Y��S�F�\�aU���{��;<��X�g��^:����QV�Ұ�&�拑�{�	��|)�J����\X�k��fH�Jz�^ܕ泃���R��� �)1��k3Ln(# �T�+b!3�Hw�h��$8�ǡŋ�G� �@�!���������+� ��W���.8=����9��/�t򬥢�|�"��(g����}G��D�����6��s�>e�B�.+Wl&���7cӥ�Qo|+�Q\ �����K�=�S^��Ӗ�
�����n\��x�F
eo2�*���N��Y���� o`�R�������N	I��bS��8Q��(z���ݷ�d�&�Ѣ�{���9j��0�>���0��2�D��[&��o��������9�<�2�4��ly��t�3�.�f�Ot��B�;k�¤:5��0N�4[Æ���x�s��*�`@�o�]��:|AE�� �KZ�_��,�z��%Pݦ���LGK娏�Yh��x%WY�U�W�<4��E���#!�e����u��A��؉y1 O�����5�E��J�`���Tgz23xT�5ܞ��\S�E�aA-�d1%�����qXBs�R�u���#�C�lݸ	��3]-tG�� ��۲���	�1$kh���%X������ `��V�K�y%D|���$��R�ena�y���p��"��w�L��'��MV��<�� A}^b5�g�y{Kz�с�E .�%5��&��+����g"d�E�P'2��kp3��
�^M�2r�RX֐��gMn�q����!-5)���j3��t�骟%m���� ����~��aE&S��Pi}��)�O^b/���(7�R�ؐ"A$7�����mA��|�;e�r��W� �e�t������,���(Jx��~g.�J�r]FRiھށN"����(R�d��y��NS���=�:��7���EW5���x@�:�Ȑ?K��?��Q���n�y�Q7n*�H��zk,�[��ʓ��R�u�Tȫ
K��
[�)$_�P׮̫�ʿ�<�m0��KAE��0��5N{��oY�Z'+5�Dg�-��8|L�2�
�#���"��
���U愤�o`���
c�JGc��չ�m�sM��V*ml�?6��T,�����X;�����/����C�W��$�P�}L�NH6�@���?Զ^�q_�{	���K�r|�	'�p��&BnW�I@e�x�{�E)�=�D��������ӫ��!��)8-A��*��FT�S�˵
��\f<+	#����A~��Gi����3 �.������o��͑Y�>K�U-�5Q��׆*j}��#����R����uA�xͿ������k�7f��;��xuH�� V���/���R-�����#��E���Zk���nx���JN�� �#���q��I�v�F��o	�C3,:�*�tK�`e�.RE�.��w~y0u!�ذ>_V�=Jә�B
��}�B�Ƚ����XI�&���A��`����C�+"'�P;�b��d���d���obW�7�]ǟ�'��hAI=;�W7���g:�����X{fҠ�W�S����ЮHVs]V�F)���bf��z�}��;'�9�r��5��M�q,Ɗ^��D�����jX�cj�%�4jꇳ�<%�9�,g���F���*�5ѩ%���~��������3;|�#YI����~g��8���ɼn�9�lCh>Ck�/��%e�+�������+��z�F��uq�{�bl�~�1�W�L���u� ^��/�+����F����!����#�p��l%~�<��,e��>�{zqbq-ţe��:'AC*�bv�	����o�Q�t,?(�G;)�������X@	� j��Vg�m�{OcR*�!&Ā��e�	=�}h?кm�P��MF�+E��*=оn=C]��?�R?֎��Ȇ]�����^��	v�It�;ɭ�ONh0_�b%�� H�@E���-��d߃ŕ$����xL�U��I3�Η�{�\ty�����'��.߷�\����pb�B���8y:j;l��ҡ��.֦��^�I�uG8A�ut�AK?�4���J0{�_;hQ�3�h=���h�<<�D�o<Q ��G�'�o�(M��� ��pE)�)��.SBM����DpQ"�@�i���{�n/���.�.$g�RXm�h��:tm���fY��Q@.�]t��2(3Ƴ�F@��'$�R��sxp�ƉLj`�:5.|g�x�ױ�X�Z{���+�/��ݫ��7��jj��n%���O�Ef�='[�7�=d�f�ǅ�eI(%�pb�xa�W���t�t(4���3I(�=h��#��U��ܺ���9�[d��Gx�HS(����ɦ�=�
H� �����Un���CB��� Chۚ�k���KطD�I�tU�&N���4{�fU���=��N�������q�6�����V�!��T_���W��C���%+�K�� ~I���� �B��*mۉ�I��y�~�ƿ�N�O�Ŵ#��=��F��p�'���6;��g��8GT"�G�qF����4��%�5�]��2�uچn���s� �3s���?����"��b�e�ya�N_�2�;�C������k�[�>�G�!~�T-��'�|WO�������+��s��s�!��b��&^*hZؙ;V�˔`��4�o�bu��i�P��4�`�~�tc��Q����{>Z�C�	�w4a� � �7���6A�Z�$�i�є�|�_Q;ЬU]\J��l��Tl���D��z2}׏���6p�����\�I{r���¼a�&b��������08�\eIVg��7�h���k���u��М G��Z�����&�J궫ږh\o�f�+�� ϛ�6p�g1�
2�/�`�d9���(��>p�w�Ac�$�q�O�]�fdt���5L�\�i"�Bߩ�u��t\��*���'P6��gm�]?ۖ�x����m�r����٭���������9#��|UΛs��ȫ�D�^�۫y�^[�c�ߌ�3����2�B�)� )-��~�����&(�F�2I�c�hy*D�h�h�������RA�<Ǿ��[�ph-	�3���;�LvS���2^�gx�X_�F?�Ղ8�3oq�(V�>�����`:�>c�/&��ALсt=��m��kYTB��2��/��-+x��]Ln(�h.������1"J�!���Иwb���[��mţ�X����oz�w"!1-琿�s�:f�i�:��LÚ��-H{�Ӷ�;��R�6���݌H���~�*;]��X�XEL��Z_�;T��cd�`����m������6��w6��Sv+��6�-N=e���;[s�m�̎b���{�	#��Q
�G�V�u���L�H
�nPa��n�n��,:��'��NT:���@��2:TZ�*;��}��7x ��g;�	�g	��ֲ$�)�]�5�nmV:��i�\��ɒ�qU?�� �_41.�kT� x�A���(������������BK֭o]��l����A�v>���7F����D"��� �@�G�	TG�|����ʹ�����97	�
Ǔ2S���-���֥���jW�4�i�z	��g��*���l��*GbvpS�wR�W��W�m���]�������|`��Wj]R[�Կ
���E<�I�U!"e��ۅ�1x:W�z�\�*��
���7}��!|D�{�O��!���fŻ�����>?�0h_7�c=A�1j��
�^/Xު�C�;W^�9O	i��i��T3�s|0,�2��G�C��5'��yY��ޡZ6maz��H8��̀���_�D�UA�;=ym 8@|*g�r:��7��~��M鑇�J:XY"�3�ԃz��ڤ�}��e�g��%M4�<�}���!n�jl{܁�Õ�E�@6�<ރ�ü['`y��JD���Mul�xjl��J7gó�-r9!������5�S��a:mif�� (agK�Z��f�B���7��/vCk��Yy��tܤu�io��=���bu����#9Tm'W6���zrTm	̀��椄M|���N!�|nB�M��G������PH�����YŸs+
��|�3Ϛ� EA�������ᢦ�$�N�@��p[
O�2"V|m_/���ڜ�馘4�f�G �f.���Gh-��j6�zZ�����������z�ӫ�|�[n��]��8�5��!��h]�+���̲FF���ҎL��x�1{;������ʡ��QNb�~���jc�,�b���삠�qb?R��,*4��F����3��
���q�=m��.��~s��8΂���q5��![�����Ϣ�h����԰8�{�&f�j�c��;ъP�[����V�q�%ص���ZI.��!x�80&�U1he���*s��D-�T�0Y!����#5�[�)��P�_�+��B2u�������B1|���?�$EZ��/�CwQ���/��G��� b������@G�§-M�B�y�1LA~ W\��O0��H���*x�����6�P@h
�ay���:�[w�t�$�~(ñM(}i�'@��D${E(��-�.wtH�J�w�rs����H������I+�.�Hv�'�����1{EXv���nHy&T���^��UƐ���R �������F�E����"��#���7�1гD�+T*n@�?��{öU&x*��C2��5�^�WE�Y��Sr�����-�����In��W�O�:)G�Q�|I�2�f�-bٍ�[�&�{�vb��:��������K#ȥ�'�:�J�>=k_S*��2 o�h���RO�^�]�F��r]��<>�N˖��	�f�a�gJ���+Ƭ^}�T���o�/ȪF#�NL"�N���{�w����m7j�q:n�H
%�OhU��jp_V�Tx�[�&F�Sˆg�+0wp�ivDe�Vlu��A>H��N	�)�$�l�qҥG�_�'� p�Lz(�ϒ0�7��/{5d�@f�٨�?�=�n���Ƞf&|�e�������.`�����B ^�T�Y��e���! ՛��-�Fb�(����L�a������_)�N�X.�	D�� ���N]��H�S�z�ǱX�9�8���{Y�jz���F��)�\;��v���_-3)�m�"�w�>T��h_R������K��
O�12�r�:�3��D���1���5"+�ׇ����~��q��XF��m�E�|�e�׭�o!�Èz`_ ���Hk���"���C���%U�,۫���9̎��]�'�����4��V;�_�:
��%KwS�H$ۏ�zD/���4�wՓ��HR�!�QǠ`I�� p=·�_����z��~�6%:K��Ь�*a~�"�D���+�L��щ�1w��9b���.UYrW_<7K��S��K�~� ��)��'�G��!�G�<�3��g�9{���,�xP+f��TL��zX�����#��o��[7�%gW�������r����r�� r 
���q,x�Y�g8���&�� �еqvaњ��ɓ��bܦ`�P_�mK��Gb�1�5�%?
i9�0�9�r��қ��R{ŀ��7z2��nHBĸ3}�1
l�و>kOw2����5rw���PW�ڴ^N�������������ܓIaJ3zI�m��7�0Py�����^�1�s
ǯ��'닱'4
�F� ��!v���=Wi6��':���<9fO����zg�4:̈́$��L�#	Y�o|U�UO��u=ӽ�+���h�tf򖿢㜝MZI�ߵ$�3R*ۓ0ؖ��� _g������Xxe�o_}�7*������C2�%p'>�R��j�#���
m(�Bse6F����bd)��7>\+�ȷYS��� 9���xJ���= SD���t�����}%�noV��&���3E����z^W� ,�2D�׎��&�� ��<-\�\@ky$D}A�}�R9���bt?���
�yrY���*.p�w�p%�$:?"N��p��q��F��lh����	���)�����|�j_�'
p�p�@������X�j�#�s��y� ��<?j#�2���ڷ2��|�5�}(><��t���{>q���r�R��	X�����l��m�;%J�=�ԗK ���~������Y�՝�}ǐ�K�n~m���z�-0N���S�E��S�����S�&�7r�Q�� ���k��b`q�Z�A�����=�RS&&C�9RpD]��>�R�O��4�%G`�
��Cz]shʗ'§�4��?�^H�Gv]TP�	ԏ��ۧA�i�O\�NClF��u{o��'�ƙL��m����γ��tT��	�\70�#�S��=G��_��Gg�R�P���B��r���p�Q:V#��yڃV�n�����5�Yt�
�����S�3���˯���:!j|'F��G�K�A<s�`|�)"^���
~dS���l+㐓0u���J���}��|��%}~<gy�`�&�n�2��*+d"��B���E��kL�2��I�`*_�%���� ێ`�w�&���ɱy���c<&�
��q��pV籔%Ju.q9-�n-Y�!x�`�Ta=����};8`$+�70�9q1�p`��3Kbq�R�˄�'��:��|�ǦD�cs��0ZB��OƹޅO�'O��9%UI���V�MiOq��<�RBx⫶~>w�.�%\gZ�O�(p�<�b7?��˱N&)<Ug=x_{ǈ�f�5g���){e���'�Ϫ������}t8Y^�#(k-�4�p�2�<�]�W�qRd@Z6�"���Q��[[��v[_DS������l#��pgaD���J��x}A�1� �@Hs�g�c�ka���[��\g��
�~P��Cϻ�Đ����w���Xx�s��Ŋ.)�!.�@dN�r,jc:��d"?X�=���w�7��ī����.'���k`��'86W �Nś���1Z:����3���ĸ^�{�yf~�ԧ�[�^{�{n�������k�ҖbK�l/�\�]�3g�Tc���D׶JoYP�O�,|w���S�����{욺�a�{H�V*j��QxTQxȕ sbړa�҅�ݹ?��e�c	a_T�� {��^�B>|O�V�m�O1������wӇ�5������.��,h[a(3'�i�-�U|>�0�a���\CMv�D���p��M��bJ��Ec�pio)�����D  E�E�㍴��#�&���U8��цk�ϳ0?�3�?&�C��8�w�f����N?�J�7�#�v�8�����1�[��� ��^E{R�M�lT�@�R�nP���pI~�>߄\*�ڗ�iasz�7�c�'��SYg��/)��pX����W�1�/מE��<8����QH"K^�yZ�l��蜅��b���{�s �/�G�[Qd�T$�[�~����)ޤpg2�!BV��q/Aq�n���ש��&�I��`��Y}8���E�h�	ױ�	�Ќ1��l���Y"Tz�p(R=��\�� �u��m��Ӕ%=�k��-}K�h��7-�`�+��ֽ�_IJr��CYWP(݊AٶF�5ӂ��0�\���l(�*)�醗 ��A�	%|�hI��-$S�YFŧ��B��&C�k�6 ����w�4��v�kY����V�ǁ$���BȢl��[�ؼ��$��]�1t_ůJ�;�����,Ae��$��)W
�z��4A��)���]�_Ol��݄񎎆W�Tg�'}k(b�������R�������t��8�,�ac֦}K��L��y��:\A�����4z��%�P���@�݆�8��u�C��z�`�q��d�C�t�1��J-k�ێ�������f8v��a֠����	�O�0@p	�y'���Q��m�*��f〧.�b�	h����"�R錐&V�l��Țh['<J��7�=j����۾��&DR�>4[M��?9%B�8�U�[owP]�7�_�tjτ2����b���m�klu$>|�L��Pa�>M��,�Y0��/��?�U��sNЎ�w���L�;�qb9ƍ5T�81Ǉ��a�� ���_[���0=ʻ-�J.���A�0�f���	LT��w���)]ZF9��|mmw�>e��hw�"�O?�[�� �f_w�q�����Θ�T�z���|�7�8,�g�B:��!�|of{2z�h�<�E�� �R��0�(/��| ��83U	J��sA�W�꣡m����I�X�!�a&�a}��4w���w�H��� qY�w��B��׊�!\$;�=4����2/�Awɯ�Y��� W��8MQg�Z]sb���T�ȗc��D
\��p�΅wĝp�2�Q�,�t�i�$OL�������L t���_�-iq�#�Q𣎓6�����IY��*B?%|p�w�E���n.�?�� -��.����(��ϵc\�W�YE$Z���J��~��}�����4Y����g3��D�y�u�G�IJ+ë����,�r���m�M+�?薉p���4,���&Z�]
��|h��;�i�̰+���elK�~���cs�Fk
N�g��i��3�d���.=c4Iئ�k�ըL��$��6(�i%�kq��!Wo"�W��ʅ=����"����y,iS0�]A�c�������N�j�)f��J���S[pc*���Ct�b��7���38c�3?���j��RLtōu�::���זrۨ?{ɑ<�Y苈�a��R�́�SFg��u0���\����r�v>z�/.����?@Z�&bA� k��ś�E�B6�x������7:���o�+� k#5��	��qq�(ĵm�q��[�`�i�9�.����_�Z�����
{����sNu�P���ːǧ�1� �{"��u:�O��� s�S����f;j����������<F2UG"�x/���^ցc���g q9,�A�v;�1�NA�=����s�=ZR���a�{�)T*��Dr���,\B����1=�5���X���5 ��R�`����(��/�|�Q*����}�\�� ��	㢩��ŤjW��
��X?�/%dz����T�l}	����^��{,�"7�fM�3���Qߣ��w�"+e�C�P�3V�sO
�N�T�{��kUH�����ש���"Za���ENɶ�L(�����{I�����O��V��;���YgJ�����""���e�bE3*��8m��9��՛�ϛKi�����Վ*����}�`!i�V�?f�-�0Y���bT_W����-t&v����ڗ��=v��q=V�u2 �(f�^\#u��3�YP�UC�-a�SU��j�W��)H�v��P'��Ȳ�qWgY`8�)pE �-����>IK�X�ŉEPI�C���i��z���$�g�e�:8�@px��~���s��H�D�e�d��f#�4m�:^�q�������>�k�n�R3��k����&�_Z;��$8��v�E�0�]1�>h!a]V?<t���,�NOQР�3�h�0y���W����@72[�o�����J����c��� ��Q[�Ȳz�G�o�|�F��1�ɠ3P��1=���&�g�jG�y7lˑ�\^l<��ȿ��-�U��C7��cCC_u0��Lv�ƺ҃S39()�FY`S�BΨ�Âj�d��W�`H|^*0N�ţ�b����M:���R��d Q�Q|�5=zR�B������WŐ��"�xt?�-�B!�(���*#
������C���yWz"$n�f��iq;��]d���U�J��x�[\�V M�<��s�o����V�a�� �Q��3'�T�l�������6Z9��P�l�\���n��/D� ���$AV��6+H[I@���Ⱦ�Z�80�6\ˋ����qСh:,�O �vK��0%igN�Wqiob��n���絏G��Э��(D������ϣ�Ŭ&K���=��ׅ�E�����=�i_�1um��9Fc�1 f xN��"���_� ����~����*�WQ����v+}Z���6�]Pt3^%=��"Y�cK�toE�Ƞt�-�K�G�<�)�M���՜�	nD�: �U��M���h�j��V'���Q�sh�Tv$Vn��c8r�y�C<�:$�9�󑓗�m-P�-l�B��^��ډԍ�"�K��:��J���jE�_���v`�ڥP{1f�W����3�#�!7��t���&H�<u��i�F��t��iԧ�&೐� ����#���H
�~����W��i �
|������Z��
�a$�~h|�fqW�B*z,��8�́*S>2�����x�9dT�D�䪘r�4R����$�\C�}�X+�c���oP��@S�)d �I�w�/�v7큺]۽D���*Wqhu:K���2��a,�WX���f����Ŵ����˱HQD�@���C
hDs��:�wh����64����壇j������.B�7vђ������+��1�D�=�f���x�Q7^�d�s1��r��ѯ��[~j�u ��
i��I��K5��A���'1;���E�OTT��= rZۉ��gW��>YW��N�(r#�)u��C�h�m6��/���S!�a��(������q �5:��&��'���yl͵�v�<���a���d��l�Ծ�toРe-5S7X�c0<�b�s#@�]-bk�2,|�q���<�*�����ى�=���Պ�����'�	;���M�)G
M0�'��+j���jDE�x>��v���X�"iw���f�D���Ƕw��g�>g&�뢡����o�6�3妞�k��4�c2GA&�b_Y$j�K���:��?(D�F$�,��ԲdbK$⛬�'EF� Q/S�$0߯sɀ��:y��`�`/g��f85�;r3lA��($:��q���IB�������+%�՛��Dx��-ܭT;G�[nC�]����|��>F��^7��Xl�� څ�|�1�zL7J.�e�N���!�(5���(u����l��đ�����)�T�&��7�S�]�Y��i(�����B���:@[K�5�#�f��kE�<軨���!�WE�g� �-�QCzOj81=�����?3�=B�)�/͉J��"���bK�R�͵Ļ]�jZ���t!Рa-�4��9�I�@gM��X�WS��HĚm�˯֗��{!�����Bww�xA`�r������]��9LU~P��Z����J����B��Q�(� SZ���!W�Wdy�a���Qh.��ݡ~��R]O^�P^v�M:I)�f���_�H������G��g1+�WU}��+�8���eZo?���l��@�5_��G���/�-֘��&D5c߻FkU�*,����H
���(�<�pw���G��_ �����A����@9�]YƤ�>p���Tb܃���+M(���8�84��ԅ2`P}^�����;l��:E�FFL�:n�HiG"�W0A_6�������^��BI�a�����Zd�-F�����I4#}��Y�C� ���+k.��ּ(��9�)0�o��Pv��rh���u"5��45q?�[����g��&��q#}"H����$��*B�y�C{�b�H2���$2'��0v0�;�!�,[������)���h^�*��߸�%���HXq>O�>65���U���a!�H�gE!�'qV=�J�>f�J�T/[$]Z�&�n����&�1��Nӆs�o���dvӛ�E�v	=���$AAMq���em|�|Agr����C�Ӵ�W�����5��}G�Mr���%""�M�iOP�U��S���Y��3��k��o�hC���CH�I)>�"��ݓmG������ ���{F:god�9>-<���C�V<ɬ|�������\XF-�'zq9��/��LZ�䊶*Ix<����[Y��D���\y:]pL�<)��C��!Z�G�)=�������@�}m�s�Ps�H����ػE
��Q�+��p�ݽ���y ڵ�m��~)�.���E$卄�B��b�07y�G��&��u��骔b�'���>���A�E"�Zuy?�ٓ>3��,	9oX��_gǵ�w�5�h,�)�x4p��Hbt�
=���EI��v�K�(���	~���E`�A��ݙ�`���N�ڃG��l�F����RY�U�F�� zEW��q�@Ю�&���&��	B����d�{1V8�(��d'(�|TH8}.i��#�>4����	2
�+�c��"����̀kX��z\4�P�����Ƴ�ү��v�)�=�Μ=�
�C�m�l�(�B��lj�M�>���r�o̝���d��r��h���6<��|����f���֛�g?��� �c:΅��{R�Z�}˅�_���"ʩ��e��n++��\XfS6J��|�Ω^�գz�C`��(�%1��Xq��m��C� ����4�Ș:��m�"�ο��bAK%)l�1*����謥�h熖́w{;����5TP����a%����]� N��-�΀!�9Ϯ����2C��ʰ���|/�B�3��LA�����&�G� �(O ���F��5��K�Dd�-��S������פr�U�w�ȥ4bܻ�����0��)��"�s�ei���lV: ���j���מ�է��+�l��V�k�{&����5u�>-�����pv0��i��u-9�%��"�fn�� S` ��Zƕ_"y������w�
�Xk�ML����S��(��bX:\��&?/��o���և�Ix��C�T	��w'����q�N�t3�D�
�doq� ʖt���~>�:�^�ź-oф��Hm��I�}ѭ��T��%����{��+DH
?4�����>������C[�m��GN̲����%n鍪��vQ�|[��ȓ1;����n�iB[����g"o�7�O�C���P?�E�Z�>�����\O\G�\^���M�*�����ڋ_fi\1[�j2�R��2�Y�z�?��� HU�jx�x��TC�|�G��/	�!�c"�5z��w���D����`�4�
���<���%��o��B���P� �J��M�����k�B2Wm�X\���IE�Q�1͙<�P7���&���o7�g^;B1�s�g�����f�9԰� �@ƴ���ʂ��G���7E�2��&&��^�g���-J����@����:+;j�XT5@�&><SdL��1c]"s��,BO�%�t�B{+=���~���{fJ���@��ٻ�F�7No�[e*���Y���?����v���}�X��|��h��P�sed)�������ə�홊G�k.y����Ĥ���k�\�M�n�S^�x���o�� p�pʾ&�����V�B�ynt�4@Z\�
�˂j ���ÖB�i�F좭0X�������Dq1P�yt/�� &"�mjw!�>`�B�}w\qD�hz�4%qO���勢�]��� ִ�ۈ�.x����^[ ߦgh�孯/��O���+�.S���Ǟq��H�E�kM�B�z]��#'�p���A���I��TÒE�J�헂��5C>�%�Ŏ@�#�_�!Y��@(�m[��L��rĽ﵈���86%s�����ݮFf[}驒j�*`�;ߐ$�9h����2%��d��>w	w�� ;�p���`����@�2���1�?�%Z�a	��#]#Z�)�ߦ�!��F�x^"�E2�xR����)@��݇ 1TF{@+�tNہ݄��vt�I�u)���B��Ͷ��<����ǟ�ïI���aRPo��8b��ZA=|p߱O_ ����6Y����г���t=s~b
#hz�8��6����'G#j�f��[<;�ʼ+��-o�����|e&K�����OBk��X�� ���o{qO{R-R�}�ŵ���i��%�,�u���x�3�7��?�v���]6�G�8u�?P` �g3��l�kT^�q��b#���%9���o+��|���-"2���̥;_�� �a��~ٮK2�0��� �m�qq�O�Lޮlȡ��{�~/ۯ ф���]~�~Q�f8{�����T���R�/�3(1k����}��_I��\p̖��rJ��@��xt�װ|&ː��!��;A��a*��Җ�[ƈ�Τ1R��+ X�y�	��p���򝨩<;��BA<��%-D�t'Q����hibt�������$���'׸��:!iC��s�p�;�ag�Uw��`���}�&�$���Q����8�d�������Y�Ѷ���KOnX%I4�=P-Ϻ���iO�����%3��K3-����Z���KIl��r��t�Q������p�! v�@��1�S���1k�M.D�����j�c�pA�
(O�i�����h"gbG�|j�WA�h�VL��gPMe^�]����di��)r�<(�[z�@4#�]���\���������:c�Z��#Ԁ��'|�āV?�ZiazO��D6�a9�F'�^;�SV�eShU�ǙXe���Z�LE�c��>�Oٳ���Ё
����n��ʂ�xt��!<3�����g��N�/�پ�'}^���(�-�R�d&��3�5!�d�<G�CM����-�C��
g6�F�VEK���5��׎�ٛ�?�b)��­%DG�1��f���}Y�˭<�� )@�F���&�~%��i&��4?i�e|����֐���d�*{�,]���[(�=�!��/?Ѧ�r�\Mϸ�P�_	��b!���n�v�)ػ:Q�My�@�ֺS\��Kc��������I�˵�����@[��vY%�U�щ� �����ϛL`���A; �7�=���6��0�����_@XW�Ŕ�M���wn х��%�+!I�_h\i�5mq�m�>��>҆�5&��O����'������&*8�^G���в+?V�T�CG��z#/{�^4K,:ʛH�ש��aF7H�m�V�||�X��)��Տl��4#�� �w&~�)���qXy�rk�Q��?kKO������!�	����T���ߢ���@�^�$#�=2�P�;���F����=�_,�E4�-s-��q���Q!O�ݸ%Z��̤֝fY�lK_Ȑ��"�����'p6Ζ?�;م�+B��?0�v��L ���o��ۍ��z� �C��tl`����T�RF��%�R�,���$��a����x	���t^�J3����Z��)���)�NQ�@�{؋۩�Lp��B���qx��D�erP�P���ԡ�x��F�����:�Zߛўʔo���C��)&@x~R��Q�����y��Lܼ��E���q�ŉ�r6��5�ɡ������W/�*��Eyj#���Fl�b�T3��n���͏7����M�A�>;�5l�Xԃ�Ix-�4tl�9dŴ,�2�/�,<��Z��q��?̴�ϱW�l�u�k\�bxu"�Ȟ�&��7j��~����nY��Nj����@|�m�92:ȩ�L��0�.�������
�/fw�E0�o�G���="�����0��&�^��qS���贑��ݿ�MM��_;+>N�1۵��MÁ"pE��Y�,�fP�o��2��������(G��".�G�-Y�$��L�߸�Ϥ9ᅨTEcWl/�4I)J�rR(�'�+�	�Xn
�9�h����@{�����vĝ�3��K����_�')hQ�ni�^���=��Via�7L���%�B��v�Sn�yEL�!HK��m.��.ؼ���g�1�%�p���w=V��2�֚��%�0F�\���gfT%1*����1��и���y�E#�/T���K�YT��%�� +��e��>�E|��qw�(!K�c��f����k^�D�J׿�+����:���͕���F����),"�������$߂k�w!�Oϰ
��:���wͺ�nɭ��Cջ?��̩vɓd��ƕl�N=�5������)Qj�"懚K��U�|~���aD_g�X�lF{�ϮI��d��>�(���a��]͓M���N�	/��R��Q�1>nL���u8f���=[6���3���|lD"]��R0m=K8X��.ؼ��&�TQ���l���"��}������/5����,����x�N/�$���v�]�������$�!��0���Yl������g�:��5\W�<��`�NXsbFJ��ߗ���?	͸��|��n]�m�	���a֒�$,x�Qw���\�iW����e�<�5-H .:kg�\�ڧ�IV9��V{gSK��d���f*�I�i�P&�F˻Q���嶐]pe��@s�f̢X�5Y���J�8�r��E����X��y$�V'o�q��������f�J1X]��ڇW%#�sk��"PUm|\���-g� Q���r�R�[=��`��Q�͓��
O�NK%ٰG>w"$fG���35��;Y�oS -�DC�,=PW�^��Ǔ3(���"2�e��3 �-�S��2_�;\�H�_	�H|�[�v���i���Nx3ϒe����ţ͞]���a�s4����'�a�X�3�����Zb�f%w�uIT
� ��Y���?�H"ܝ��":Hݨ���~e�--%�FR�>4i�
�;!�c5R��Y����t�/�Q<�����F��bg���b��u��F�u�)]�E����s�[�~�=Ov|1�?�~6�g�|���;{��N�Ma2�t6r�Z\;�k���=���
��Y�#�Os�-Ծc)�7�<�oQ�r���I��tXl޴�D�P�M�J�2��쾿��nW�X�.�ӥ��l������D�la�?{♙�jjAN��8fh��͵�9T6A�8�ث ���	=��?!Εg`/�H��J�l9�8����@� ]O���5(��EG_��1����Ĕu5�)0Ы��˳���HW��-��}�X�ۃ5�>) ��=�5é��P��fӭC�9GS�=������+K�4��Ӗ�x���Um)a��D[�ߛͰ2lC���0o�k~�lb$;W�#EF� �O�E��.�:��8\��jk7�~�6�,�i���4%\ny��!7H�`*�f�K���*��C�P�1��F��,�V�k>Icb��������mzT O:<�7߈T'w�-�7v���W�M]�. �Yr���rh�LF�*v���G�����s@��X�%?�IA�`�n��!�_�5�D�Qt0�	��c�y���'�/�3�3%�5��	M5;�BI��k�7�c_Ta����W"#��zcȐxg]4��C����;�����Z֤�S]����!��{�8����T�{�1����K�h��ǜ�n4V�8*�����"���G�C�����F��ƣ'B��H$�M-��5�|r43�<�F�1X~�+g�"�9U��8�)褞�ʉ-f)����G��W��uߋ)a�1�;Y�pS�]P >q3�k[r�B)&��cğ��5��I'�@
��Ta�!�K�����^��J�>ʩ�.�F�_��BN{��2���l�KYg���NE��M��.%7�Y5.���<��?�����]Lϥj+a�������W.
;��L���i�n@���o��H���ƴxE�M���j���{8dz|�SPU�2��`��4
�ku�7���1�k��q��O��>��w�x�S� *(��l�	��=<>o|�S!F����A�7�����	�k�%�]��Z<)�3laX�At^nCЉ�I�K�����ѨL���K��x�ݙ�?��+&��m�7D��J�����#�ﴪ���*�Ȁ���|4v�7=.����"LU8��$F�:p8�<G#�Q����l���Ҙ�e��Mţ��3��@�l�D�6��1�T����(��o��1��ŭ������a�������oz���.J�?�A����M��H��!��-]ko�m�Nθ�ފC߲����,�.�S���!
�6;��C��|�ٞ2�0��v`�q���N�ro:�dֳ�C51T��?���n�Pȭ�������X�N�`y�6Ja����N�S��U<�:{?=˶X��E[��X�W��v��%�.ێ�߰ٱ����~[�a��6!���?�=L
}���K�f@�hm�[F�yA9�����@걷M�����1�Y)���2Kq@��Yl�~bSg�@Q�~�fW)#jE|��Af��!�P�[��Q�mq��$BO�T �/cd˶e�v�#�?{��5��Q6���a�!E�k��ī|��@ꝵI�;S� 8^�+qǋ�n��wTÙ_�Q@:��Ҿ|� jW�T��D��N�L~��.^�Y�@�w��hңW��n��9!�wB��5�D�w|��7oG)�R������&�%�S�<F��R����E�:�D�B�t+{76�xq"��C#ğ��-���la�ף�Ӓ��m�^�dP�`�Ms��֧&�b(��_5�"F
��gj�������1�?��+?���:<��P&���u��'�B��f����}����]��R�؂��C����x�k1��A��6.�ID��|Y��EX��i�4������"U�u4&��h�H *�"v���x�\C�E���2�ٜ�lj�m�kb��� �Z�ZRo��C�Ћ�����%rZ��M�.o�YV�n9� g	�5��.��go��?�����h������b�M�mnR�'�2'�'F|Xs�E	�cߥG
��+FI溜��=����$��2��H�S��D�QC.�v  � ��)g6��7���<��'#!���k�i�Z(��,m���o�h�p.7���g,V~��B�9:t�J/O�T�H$H�a�ݞ��A��ClfX��j�j��H|w�6�:E7��:�n�w���*}��P�.�Ӛ�<�w�î����?i�s�6����eKJ��J���)0����M�[W�3&[�1����+���L��9J�V�<]��Bo�| &0�^��k� �,'��n���Q�4��@���)�5F{��vj+�oSS�����'	�uWB�x�s�?�o�ԃ�$�!�̇��@��C���F�<�����[5B���L̙`�Z��F�J��ȹ�ͮ�6�e��T�r
�	���l�2n�"90#��?���K�3��4a��,K+,8�ٻVr�٣(��Z�Yx��"��h�`�2t��i>N�.=ȵ�Ta҃������~�
JJ�g�@�ޑ��.w�?Pʥ6OA�\!��iS�4���@�Tw:�U��(zѝ�Z`�!Zm�򽼡��1Y�L�ww}��:e��#wp�Ӌڞ����g�����d<dH�-���)���i|����xL�D4	%����*^\jT{Y6��1�6"E��*h�nu�K�5�i�|�[��.#��Π��a�	і7�����1a��g�����u��Yٵ3�J�V�x�`D��d��z�tHE�0ޕ�2��0��R�]�5���{���p@�|�\6M1�R�}����.^���3��3o*{-�´�3����&م|���b̦��w�	��z��7��En�6��jo&�ſf�b�y�S{�!�*�.zc�$;�d�E9:oW��jM�3�(@��0�Q`���J�B��1����&�0�x��K�\��D�į]��A��� �2����y�nF��9۲]�M�<G��4����O>1��0�j�u��Y�U�{����Q��M��g	���i�F���h��Jo)qW�z��H>вlI& �'R𝇕?����	U�:�^_`��O���V�Y�ekc����.S���P����t}�2����k�Z� ��|m�Q�Ll��kQ.<����~��l����,o�g��o�4�
�A[����j�w6�BN�k\Ξ��Uהe[uLd��z�.>��� ,�H��>�2��T��G��W�.Z:�����񚡟'%��n��.��X�o���P2��H�M⭩���=���n�%��N��ˊt)i'b�$E�	(�.1�3#�}P�X�doSC��7������1e�ϗ�;���������L���3K�Vr�'�=�<I ����6�"�i�>��X�~��Y	[�y�����bs�d~G���7�����1F���pTͣ?�����Hg|BL���p9k⚴@�x�[�B�0�gd�8��¦�;MǺ\��0�t�ʭFs�9� 4F���")���x��-FS��.�����ڋ�ȫk�����.B�E{�����#uqO�/�'�k$m|,t)�FWpG	�%��c1ڃ4~� �g)v�+���i�.�ģ������%Mf��×�����"B�eõe����X�6�w��f�~U"xյ�G�ȼ&������j�%�#*K+Z'/��vj���.���K���==��JA4�G9E0�Z��%�A�Ji�Rnt�_���
��݌����6�Դ�x%S��i���0�K-���:��83#��r���n��BS�,�}]n��#�I~��O�z�Q�zߠBR2�P��j�]��*s�G��������*M�1X������Z��H��l�~'2%���"�� ���[���0N?�"�]�Kh�Pwuu�/'��<��:�%���m &�m<5�F)˟;�-�&*=��6��n(b�1��r6U� p�īx�3����{�6�`�Ю��A��6�UO����y�� �@O�FO]nlvަ�H���LaIT���ݒJ�z*dV/*�Ug=Hv�'�dq;O�d��¨J����&��m�2���4�I0��蒾j?#p6A����ʯD�#��@��E߳C�q��9Ca�.��PC�Q�O10�&M����ƈTg���:ax}7P">]��׏�b�#$ǧ���ʖ�(��/���0'�	 �r�0g`Zn7W�������&�}<�JDf�>E�)7�(I  e�&�Q���ϧbc�=�6�ңs(Z?�@���Щ��4bx6H��d�-���q�-��ҳ��i���4�s��s��n�#��'��?#z��:j=�m�<�*7<R��2���
���/���-�+e�
�����rfg�Y��9mX!��+o����3�H�Q5H�_a�~B��@���:b*���9U�E�uW��#S�� �����Y&�/�q��ֻ�,9\mO�'`��dY�������r��hx��<ݓ�5z�\�#��J������(X82[#�)W>��|{��3��o#�-)�$ЛY��T�ҡ�t�c��Jr�'��~�nJ��$���8d$����Lf�gz�0a��_s���� �݁.��&t�z�.#Ȕ��5�]�]��<e� +`;����!�iFt*M�@�IeF���Pv�����m�K���Z=��ё!!,�O��� ʧa�}S���ȉ8wk��$�+���#xxta�X�8�3H�+��[l��(}���<)��	�%���?���|3�dư^���^��w�&O[���(?�Hݩ<���+h��� a�|�i6��Ɏ�Fվ��s��O�+���.^����qG����v'�6�Z�����d���]ޯ����.!�;�1���_�Β�-0F�Gb�R8��Sz~T���)R����֎�@u�lx���\�i�g��f�S(E�)ܩW���5?�?��k-���u���d���/�?�9(���8� +�/-c_l
IܿNǡe%�|z����G��p�j�+-ڧ���<}�Eb�i�xЄ?	A��pƐRC��!Dn����Z�ps&uJ蛣"�v�4�`ɇ
hr�b��5	Fe��\}��$��-�̎�RX�2�b�8
���lM�dI5_)zzꉗ����y����H���\���C3ϖ�t.������S\�36�mR�\.*�����eq9����C�_��+30��W*GVqՓ��-����q�m���?޺p�W �'��#�;8��xļF���j��r�Rԅl��՘��X�X�n�����xS�xg�z� M�q�*�7�e�[�Mg#O@�}�S$�-S�]���y��:KD(s�~�a��¬.�3����Ӈw.Bo��)t(˷�̈́7
HN��iD�3�c�)ASu�G@$p/��0��fsm����v��q���8a�mZm��1�O����Wm���o�,������XP�!4���o~�E ژL1.��RxN`�s,���eHoC$H��[���k�΃�G��CHV����;��m=���C==�x�赂2cM+6�CTe���� h�D�l�K�n�L
��6�]R���u(��> �����sX�,������8UxY��v�#�g�V��3H ���6�ɕb�n������w�F���W�?������ȕ,�2����Ю/��aO�jyI�S����hl�X���fF4�o%7��m�7��N�N���3�&���f�!:��2&n�\��CJ�co�����#��Y;
�x ����A��S/W��M?�~|B"E�#���'����ב�5�`fVe���3[������ �S�A�����p����n0�����Gb�F�}J�$�/�l�w'��f��">x��H��� ��d������������d]n�bu��Y�^��}��Q5(�x�8�Y����o)��B}��La��9��j|����D�����q?cM):�����/AHu�Bm��]��<�Y�\���N2�F��>�Ң��@����w��ANl	��ޓ�]���tUH0S3A�\(^�St�����Pb��d1�u_{0��S�W��")����X�rEgI���M�#�u�n�t�{�$�{�&mOKc��q�-�,��|5%S��GC)��ԃ~d.ȹ%�+�M�X��e�1��8�g�[�4R~f?l/���� �� kܝ��L�G�,��N��Y���E���e�����x7_�����Y�P��ܨ�	�EҖ'g1]�7�B\V�qt*� ���
�FS#���o#�H�FH-�y��i�s�-j« ��u�;��*рhP�7�Ruq�\Y}�����΋�7D�,���Cȴ���pHX㢘�봬Q|S�a���8��ǚ��Ł�p�к �F�.]��AC�Q�ٯ��@��x`2_9����C�PE5��y�($��Wj������Ɠ��-.�D�6b
C>���ח�OthF�*
%u
�|���w^4b ׎��[=���FZ��X���T��ԗ�픱	����;�!���S_�tS+Tb(���Y�-��������o�9.���� =lc��;�<��,nWa��/�s��Kg9��� ]�̑n�r�́��"fTB(b&�����,5�n�v>v�59�#i��\z`�2ʿ3��8a�64@�B=�t�(��7~s�0v�D8��8��=� �3+	 �sb?���3�5�WSF�QLᮀ��3U4�vď(�g#�PD���.0Tеr��ٌ�d�A9K?�	��	@��ކ�?탎�n-	b��*~�r���42��oF�	�P�*�S."�%����� K`m{�Ƨ$IX�-�ǳ��G��l/�d�e���Ug9u���C�t�#�Xt;� ŏ�J��ot0BTqaho��&Ӗ]�I芊�{yQ*�ɹ%/hv9UA�����X����2� �h�.�ȹ����V{����jB`ݬ��p�.�+o�(�xҜ
���F��E_;>���Aґs�f����] �!�ec_ʿ�s���5G?آ� gX)w�Њ����E�� A3}��E�^@x������4?�<�w���)��vA&�t�HT����ym�՚IM2k�,�IW���Í%^0��{��$��?��@�7,s���mzSo}|Ķ̜g����E�ӗed
��٣T�Q_�G�����$-FeH���,knԡv��fB��3�����T�v[�R�����:��h�n��_�ߚ��
���=J�N_8�i�[gR��V���*$�c���ʧ�$���C <n�6H��-��ׁ8N�RF?=z�>�[$^dn���DP�J��?������Aӵ��+7�@�K��i�f�	�j������^Ul�� ��56K@�)�I�ч�5w�@^*����E����=��#�pq�a��81�ֱ18���><��޶��������#F�g`�^u���"��b ����>�8����F\�[伏r(�� �;��S�gf�y�Mo�������k�"�P�eЫ���C]'�[��lT�$����F��ׅ�+��O���6���hO��{eMa%�hB��h�{����(�
�K�B���Ssi���kO����@�M���J���4��hꊐ3���#�iT��X���-,�  �UW�|y�X��T�ў�Wt�Q�i��, �O���3��M�9�:dO�E�1��z���