��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X������r��#@�/�����4�p5���4;Od��N��r�I#��7h��$�(��?�g:�ZGY�bӍ��0Yzb0o �Β��A���p�6� �����4���eb	 ���5��G��r>��T�CF2cΎ���/�wb�!�~��R������� �1,]�z��q[ }F(V)r�P��X�~nP{o��\��L�o�'���8' r+0\>(z��;k����C�� �u���PE� �\��B��R�3cؑxe�1�S���(Z�ٕ'�[��\���u�K�?��N��ϙ@3�I�τvl�����i0<�<|%,_1�R����^�jsZ�>�~�V�ߕG��ųn��Ҋ��	]k��8 ��,�����r���C��iHJ�>h���_T`lWZ�+�u��E윖՟g$��&RO�l=��V�تPS���;*��O�����<�U�*|m�/�Gϓ����m���4���xH�Y9��E�	�p�|��6�lȴ������W6���!H�]	q�@d��ڿ�]0*�����i3�⚕o׻�=���� y$�L1��ѭ��iM�����3:��~ؤ�`�:�-�x�B�˚���@Mu0��X5�;�v�B�v�f}ԹԂ���c�>�ނ�eM��gǓ�U1<��J�������r���!���*v�*.~e�A��+Nx��[d�����u^�]F��`m�DN��hN�:?��j>���ʭ�nBtXڧč���/|�ƨ�E�����A8!˕��Yn�h���褹�H�So�@��r�a\���e��L"���r	�9�x.j�suh��W P�%�	��јJ��%'bHý�6R�i����.Ui6V_���7��xdj��b�b?�$"}�����7�L�=Pui]�#����F��n��լ�u�.h!4�ڈ ����H&�2�c���+�$W��S��9��d�u�Y��X�,~�Η����գ�_J�A�&rJ�&��3��_�wȢ g�N��6��{����W�+
h?Gd�0F�{%�v$c
����W��K����fh\*�b�:j��l���WՌu�4����$k�ρS�6L��u!E����28�a*�����*�����e 8��}B'ߡ4Lय़����b���Ʋ\Mk-e�L�8!������ɽR�j��R�_ļ�G&9��ON @C�W4}1�-�� �M��U���O9���+C�d�����5�RR�}ֹX}t_�VTM^�G��x����w�;��¨�VӾ=�o�a��H	B�����M7�ڢ�W��*�9���+�)#d��0lO�O����b��7�"���^�(V�ւ��f���7�K�W�C�?Q�]^��Wܗl1��W���f�^��&�1�b�Ȫ%���F���{�B(�T���Y���!�N��f��4b�o�n!�t����6��3����	��v&ct����V�kA�*��9��*�2t��n#�-��	�C�͖⊪+wٰv^��V�j^s\��4���WP�d^�=��
��u0�d#��4Y�����0��h� f��ǚ�J��yO!�N���EŹ �Y�v��<���e����t�1����m;�}�CP��{.�a]���B��pY�&$���GlNtq����Kq�����w�%c����1�
�,��Z`��TJ�`����é�.�Kt��ҧ�����H~:L���.]��R]	���7��J����~�nc��Ưkh��Gңښm&L��SN;��W�)���zT�P�M�_���ok�n�Б*(?Z��&��HǍ��l%e��O9�N����z��F�����`e�	��A5}���_�q8��Ⱥ��1�l�Pd���镲�+� ������߹��ם� �8�����PiN�r�O�M���p��nv>hTn��Y�(�dD"b����Gd���0U/��-i�����V?�����$��-i�
\{\(#���]pǯ�mS"��_��H+8�Q��"�߲�:��Ts�F�f��Ȏ��}5Vn:�0BwJ�(U��N��x�B�aЖ^le���r�QM��.9����(3��H�l�__�{q]�������U<?F���-��`c B�9�(,�?�oɩY��|�K��j<&�l�@QDv0�.zd�tn�������ǜ��y�Ζ!A8hEL
wj��ήSr�&z�5
@)IԠ�F
b9�Ynyc��&O�/2�So�ԧ^�{t�/ou���;x�����)��$���Ra6	T��@���A`��x��w�>K�A��j�5��+e�л�G�=�������'l%��
���"��c����j�	�_溞n驶�<�������t�����`6 �T/މ��H�:̡j��LڀȐ���T������$}@���'U����My1F�v���L�m��c�x$v�L}yPs�q��3m^v�@�8��Y���n�coa��ZY��6]�`�Ӹ
�`3N��K�dZ~�yT���e�?�d=X���2U�hX4��*b�=��?9/OB��͚+���T�TP'�ֆ�� �Xu�����u-���C.�F
�xT��Vv�)�~27�V�� ��O
�&~$cja��:� c���I�j�)5_��0��E��T�(��:���l<����b�a���U��<m��	�.��+���v����cf���A.87��Ӎ�[�c��߇���/��H�	!|����A�~�����{nv�[L���g��\vw�KS�F|��S�6`-�m&�EP18��j�t�^�p�v:`��1X�_��h\� d�������r,��������H���B��E��N�����yB�>���[�d��ٝ�E_ ���5��(ER ��m�0�]54���k��@�}��X5vҘ@ɨ�7{�����g6V	�8E���ٍ��Z������ہW��D��r����Mw�ӛ����d:#I��Q>X���2X�[3)yGe�����h.���.�f�lz�t��+��& l=ש������X�>��Z�e;�O��
Ƙ���#���m�N���܉���\EIdtF�q2ZU<�<Mx�����J�M$*ĝ��*�&�Z�+���_���z�V�%VIX�H:�����g S!�Z���2Xɻ�Fw�zg�f�ǫ}R�#.	^�(E9�Bke�m0�t+��	�>�0yG��G�ߊ�X=�Ӝ�&GD��<���T�u`�퀎����oI�H�fy6�chD5Mi��ޓ�bAu�<�4���z��s���*����:a: ~需UP�{'6�]��H�"���"B�T3ҼBl����J���'�;��U��2�6�!�ƴr�%�����v��a�~����i�z.+�bnr��l����]CdTz����]�Mg1Y^����خKa<��4��ٻ� #v�^���o��ۼ������"	�w7[�ﾁ���z���"���0,֝�|_(��Y1�T�ζ�<��in�5TڮS>.�pØ7B` 6#<��.�$�]B�<C���OřI���n�T G���^K�?�ٺX�����]�ku0x�)�7n۟AhR���Yxဌ�1�8��B�W���z���\7T+z"�y�G�8�����dd��T���5��Q(�`5�Iꡄ��`�G�"$+  �9D5F���� ��AuHg�d�TS�S)E�0c���8�0˂���u�g��K�����ט������s2�R̬�Yv]�+2AY�!sk����6��_^��!�/�"X��e�k׏��:���:�K��S���#O9�����n�H�W)�J�k�|&�>~dC�����MS�T��5�������h���)��^��M~Y0�E���$�d��+��+U���Qa���z#�P	b �M���|��T�`�5ٿ����-~�R9�m��˔�6{rQ�[&iΩg�^��8�:U,4���8x��*��Ba�k�
M��/�G]�'w���$3�>ߋ�k�24��w����l&��><�-�҈�T�|�֪Y'�(������-�W�9����ҝ �i�����Gr�?���.���ةlcFKs��8�b�5L� �v����׮GH�k'H�T�� �����i����j�����g���e _�s��9�<����,��S���| /At7����!9g���H\�pH6
n�`0�9 �Pd4p{�*�%N�J�6�]|�*��P�����d8{���k1�e��7�������^b��؃�N��SC��ZU4tQ#��_�2���� d`U-�Y�{\�=Ln�W� C�*欂��;��ˈC.��s��@��7�6&Ex���ሧ.�+�u�������ݩ� �@��(.<��fG��6�f��#X>�s�j�z&-��n�f�)MMf���;V��X���)��1�d���\eSqS�`���SF�e{���{rz��$�i�a*��G�X?@p#�U-�u�󖬩K���`��L���wq����XG3-���%��~����vo�l�<.�}��0g�oʛ���a��Ф��x�'�9�N����Ig������* ���Te9{~1��t'�1St��ju�kz��^똠DoC�Z������L���F���W��D� ��c��j�����=��k!-������4�=��}�"2hVw��w��[W��z�M�F�ȁ/ 6���[�p�0 �v�r�C��,�[59��>��<(`�8�w��d�F@��+Y��
E��z��W�����fq9�|��U����~P��8tO"��)�\����e�'F�K��"S`�Se,o&��*��v� ����1��BR�F�Ν*dyb�5><^������-�ݭ����p���cY��&@�[��$3кb�_^���g��9�[�I��e@.�s�ò��=*�=��o���־"��p���ܡ�&u>�G�h��Vp�(P���(�8.�n�j3C�Ι,�@�	l���k7�Z��dD��3��)����ջ��/�mU���\��;{a�mx����Wr}+���6ĸ2�?���,��)��_[��$e�L���v[P1��6J-�J���k+��4��{��q�m�:k��8J	����։���gtM{��{��P�>�K���	�����?��,�j�2b�۳{2�[Z��l�ij�m��!�� �e��"<�
�{g<�Ew��EULG�!��mX`:C9��
]tJ�'_�K�7Z�suU������_��6����}�D����~P.���BN�fs�a�եlĸ&@
s������43E=��2�����ے�ȟ�]��nd�}�MI�v��2/C�&�B�G�B]�OVƑD���)��A��i� P��M*u�����k��I�+o/��e�87˄�;'�dl�n���X��P5@�%�2�y�]C?X �� 5y����1!��%��gY���e�k>ζ좡)�pC\C��H"�󖳅�$�-��<�\�t`f�(�q@���Й�Y�p7�y�F��lY͆�O��$���ۧ���_`͋դă6�(�ط����W�Tu?�Ġ�g���K�"�
����hC�.7i��J�WP2�i�D*���-W���ע�O��T~��Jy�ʻ��x�r�T�䶬�^�3�}�
�����v���p����n�s�s��+�vkP��0��Ѕۙ�"�^����*bW+�1��x���(��~h����t]#@�7�f�~6��"�a&'٥��q)�1p_~��!|��ܘ��G�xM��Aǒ$��]t;�`�\t���6��s�w��d�9��-��~�:U��T�ѱ���$�I%����c�·:���Uf-s�����zK�
E���̥�y�u�db��N��~I%�Q�f�%o�ߤ�Q��IDKs
�t�z������I���x��jp��=�ǀ
~��$�*aFR/�f9[,H��~A�'27�u��S����CK�x�y"�ed���mZ% �;8�љ�_w�4ާ���+��A�fUd� �t�#B����C�h�B��6E�1#-�X,g���4�(L�'�-�V��^$�+,@��:"��ǲd���;Xi��;��ݩ�'#;������ϩ����p ���u��� fy��=�#�N��<���	����`t�$�/��+7!�-֩��ڮ���J��S}zn��vq�Nh8ٲ�6�5��L|Q����Y��9nzM��^ɨ�!���f�r�8�͠oe�Y��JlY0�`j��e[a`eQeT�*>�c!昆h �,��hD����h�X���)�Mmo�,e���I[�����脻Bb#�|��<�3��3/�).�]�� 16^�8(� ��ƩS�y��ЉZ��2a-*�{44��u���e��z+�_3}�r����.���*���t��Ħ׬a�Z�]��R��L,�x���|afٞ{�BO/��Q���Z�����e����&z3O�"[���<�;z�������a��a~)}ZE-p���pS.)�ӥ+�p��fz�E�F��E��\�p�<����M�]�S}����5Ao���jԐⱈKѝ6��8�j,](�R����&�l�yܜ�cC�]��N-�7%	�ˎ�ֲ�t��V��]�Q_��]`�%د+�����o��s\�-��j2���q#����pO�'�}Z\j}Z#Q���S��ҝ��߻M}�`h�:�̑$>-��z�m)�QQ��d�0{�D{�e#�8�8䲤�0A�5-�P4�L�pU�U\g�֤@Fs&����H��"m��1��#3Ҍ~�0D�}�^f��B*�A���nx�Y�g�3�^̚ث3Ƈ,7�Z��G0�M��1n�♑�:�!�<(
�1jJ���x/��Uل/x��
�`*6ҰI����V�n7a�j��.p\�]�����	�C����3e{��,[�+�@<FW�Ǘ��<7鸌#Nf!�s�ۙT_��ނ������J\���nFn�yI�gp�o�4l�s�>J{C�S��$LW��G��T��we����_?;}{��H.�\s��J�4��<��x�D��A�[��(qT�Q�J��M Rd#!�>m���,�'�����<���G��.�C���p~0|��1��-&��k�B[3B�V�9j���ߦ����ΨB�?�f�y6���:��ـ�cG�bgK��&d�aF�h���\��#��M�H�l���#���L_�4#��d�4q�H��)��,�yo�c�����[�F�"̌��,�+�%א�\e��n�h�d�0��K���ya���A����Q���E~О����[n(�ꦨ��0�����ٻ�-�a"�s�	�]���m�.��EC�$��n��k��$�b������Б�'��(��o�'7We���}l Ꝕ=\�'�u�uë���QQK��pd�H�J�P��~��ms�ct�2�i�{���'�VB��9�r�	�g<�+9xV���j���1�V�o�9�,3����P�hm�Y��'�ₑn���	��/�ٵ��[�v-1�`a��u0xl�=U�P��/��XQWFlة�z���E�Q�n�eqx+.�=�Y�3Ku���\R�E�G�9��O��g�+�C����1�]��.AL��y(���⽱y:����M*��+b>xH�YU(�#iт��Qt��A������r�t��|�� �0��
�Z�̓M^"H��W��#L���UC_*�[H�tE^��� �wK#�N����ˆS��db:��3�@��J �=�x��E�˟S��S.���`}�^ .���qێ^[�����k�8n�2G(ŰҥI��a�������"騜�r"�GK/,�Ij�y*,��4=&N9���!�y�����d��ŧ���1c��`SC��D��0v�
N^��V�n(�}6FR{�f�}����Q���X�  mK�҂���<8�Zy'R�ך�B��uɬP�a����3�ʹR	���+�=O��y�f-�kO����ن���{9v<�U7� �M�wL�xR�A#v�e�\_Z���� �kp�G���
9�Y-Ĉ�|+ڱ[�=����/����������� pn5)K��^}.34��fX�߼3�j��iS�n�tHEʥX�����H-���������s�u�r0"�9�����.���;#f��ޮ�8*����߈ߓ��EH���@��}WR�T�,I*9M+�|�!���T���'��Y�a��5��[�)b��<��d$�!����dU�� '�#Q�J�]����9��-���cj�ol:7q�����Etbs9��R���L�&�O�m�udkN[|1h�)'C3�]R,ߧ{���C3��h���BoJ����|}ߘ#�S�kUN���P�i�S���S�a����x�^Վ3-hi4�����	��R3�H
���M�3�hk��h��9�sD$�5�Z�q��/�Th��9���SBCJ������.�[j?�/����آ�����zZ�-1�l,����!�X���A�����g�.�>�`!?_�El�-*���R����B�]��x���^"&:����q9rGS��]_4+���v�ֈg{�����7�3<�b>�u�w�@��oK�|l̽� ���)g`���XJ�;�b��[�k�$ǇH��%��EPԭ̕
���	����Z_xek(���W�k�V�y����x^Oν��|3�p�~�Cj*Mq�	y�߃s�"�=07HzQn'�>�s�LC��-��Tq1�u1T@�xS.H޹��Z�iY��b�,���0$-�9
F*%���#�]\�sUK^�N1�O\B8��K���
a��a?A|$ڸ�[?�\疞�nȺ#��]K��%B扤85>�)�"L��`G
�(p�3%@��fbk`�Hb���`�l���T%艶�<F�����8��,v�k�Tg��ࡱ�/Δ�BÁ[
t�3�ڻ�Hd���ur S��r�n[ji��s�\X�FG/K��x]�&drik,�ߒ%���o�D���{��Jx����/Vލ��'^��Q� �*ia|����#������������ �m4��ʍ��2 }$���`Q(���7)R�� 	��s��q�s ��P��]/�����hʲx[1C�S |
��<ز��l����=
��^��nuF����SqSS��hc�@i�ih�QyՂ��d�^k����P�)*�Ij[��KJ��ƥ!�4���Es�4�o�_���9o�{tv��В#Vp��EA�t���҂�ai��A��?�p6Xi*�v�݈&�ưU*��E���3'�V�J$�� �@N�Y��跂;�	P��?o�k�I��'���妙�����-�B�ůz*��&�'c9�lp/�s9 셧�}���2�x���������	��]�`0t�{zt3�����g�ը�vf��o��
�ئP�G��NqEcS�k�������2�I���"UGUS�$v�W�5!�<�k]�*���߉X;���w2�T����h]U��Y�x�mAx E	�RL`���C�	mO�~;i�Q;W�Q�����k,x�2��M�<K�[�����W�i��~�h���zs���=���ԛU�y��>�['ű�ŭ^R �J�B&�qA��;�"K���P-�3�WAe�o���}K��'^*���VV�!LT �5�T:�U<��%��<�U�4��{pS�y��k�I��J�O|m�D�����F���|���w���]fH����p���m��v�ÿ������q!PMS��rXG����4q8�gIǶ��a��!���:E :&k���"6�ț*$u��5���)G��[�,� X*l�$i��@B\\Ps������4�$C��� 
��`��k;���K�Zⓟݶ�y��"�|��}�jۊ�悼������ĺ2	(��=���Mղ�m��k�&X����-T�N�G�@IQ���m�����Y�񸺓�9K�(x"���u�z(q���I�H�Z*?�ܷ�vEoּDB�#Ƀmf,*�=��*:'<躶O4�R����� |�C�Nb��g�Ǧ��k6�u��*�F��U�S�a�՗Hk��^�M����q-���c	�gmA�>�~�-�D�|H:t����`7��*�f85�o�r7I��$���X��?_>�8!M!YkA\+��hN@�/	��Ԙrw�B�gj<�`-��[�֎N��+�d�Y'��Ђ���ú��}���|���Mb{�e����w�����03l�j��c�Ŷ�	&J�]N�����<_�~�"7Sng^���5���Wwk�����|�'�����9�{����Jy��u�S�Q�2y��y1�$V��̃�ab���~�#ת2����_K�w�0z2��<S3�#�Z��73/��ȷ�<_J�͊����.�����yj���� ��Y��y\�xS��]���7e\n�0��؍� �zDݽRⓧt�hX76��@	�T�|]C��Ax�CH3�ư�!z���c�g>��.�R9�Mu���џ`�����ц��Ʀ��",&D�ko��D�Zo4��ƄCQw�����&�|@�%`/PN���0��w}U�e�����9����7�9�j�9Є�whxl���P���#S^�tw��I��(ΐ9�O��p�7XS��y"�~$pP't�+�������\W�J̀��?U~������3xC�B���X�j$�B�e��� �"%��"I��;2 ]�����د���^.�1��ݠAuik�z
���=P�<=��33)�� Ȍ�#������Q.�r�Sz�������)G'�G���*��;(
F���b#�%˾��1$b;K:�1�6�V�9��>Q��&������R�H�����/�)���5�"^�{��������J����D��e�æ3�l���Jb�j�!���Az>vb �����8��$��{z����S��$��\,��G��B��ڼ���јz�^�tr���ٮťg���O0D����̒�,��M�^:��.�V ֢r��E������<łJ?�y�d�ywy�lJ	|�����U�x�-� ��m2��X?"���b���(��O�L��J�p@�v�qC��\������j�H��f���Ǜ������wp_�^Ɓ���Jj���wCgH���Q�{�b�Gf�~���(yP˞J���g��x���ҽTp�lR�~jp�Zp�;�4�7S��-hB�N�����>6H'�!������5O�67��m}��~�����;L+�<�H�����!��+G���0��K~�7�H�[��h��sM57om�y�0���l��6t��g���F�糈Ru~��5���JJF�7LZ� �̯�w��l9��B�Ĺ�Ț��,ߡ΀���;"줭�}���T[��Ѹ�g��U<�$��-��O��D��I�l���j*B�V<L`��*fI�M"Xe�
;�$�)�N%�Dx�_�Yc�/)8&����l�r�<7�D���4�i����{ު��-�}-�r$X���}���UۯH;fn�_1��5S�{�e��G��#N&�z�ʨ�d"��-�ك��9{LJ��jc>`�w�"���j�=�m�J���я�U�E˘��@��u�Z[J����{���y�-�.����M��t�>(���I�]��\#�ʨ��ub���kf;ft}��R�\���Hcb񟩔�PG�%|��v>��z>�R����C�ʐV�2�6�z1��yj�IN�jH�r���e9�����{�A�6���(]�)SD}�?<�m2��h����u�C�r���OmW/�
�%�-�5� � Ό&Mք��FW\�f
H�*<�x� ӷ��E.��i6��b�v���W��>������Y��%�P(7e��X|�ʱ)�Z�H����
@��Dn�����ϪkD8��U,��ΉB��� ����_ߋԤ5����4.����B�pwafk�4���Fz!m����Rw2�R�Ƽ]�OF���0�u�.���v	�n�����`�"�E��\�*7��n@]wc��堾M$����Bp�"Ip��<�eI�:x��c���N�9\Rv�&��O�q+!M\A�
�������'l�D�}�E9,a�ˢ	�y�܎��zI4�j�3�o�(V#�{)����r�D1d�m���r�?�?2��}�=�q͖}��5k�u&�Q�S��O��=�T�i�Z��{�綍�R��E�wV�2�S%�P�Fv׸�>B2J�Bh���C��/%�ռ	@��Ѻ-���87p3ޚ�P���HA`,Gx�EA�h�MD�ߍw�J�*���X�L`,��v��z1�V^�"�%h\Z���}]��،�&X�iXZ	9����:l���w�����]M��h���y�[D��$�օԸ|��z�i)� �֞����PO����.m�[�E�U�r&�S�\X�����E0��@�O�����D��d�x��tA����,���ЍH�%A�{Rz�a�O�w�Q�,
�b(8��1?1vN���yS�\ϱ۞P��OY5�K?u`���U����p菘 ��mx���bX�!8��� Ò+X� �*
~ݬI5�5W�i���3��J}'fP��dC�9�g���o���&����'�cb����
T
I����^���#i�w@�[<�6-���P���Q�jz��1�?�8�w���_Z)V���a�o��W�2�i_�lA��d����c��g�z=����V��X�c��X������d����_2ϦZ�ԗ�� y��,���z��)�%�Ѓ��y�2�f~
��W���/S��f�K��%�!H�i��)R[}���3,X�va�n����|8��D��k��A�#�bZ�˗�6��֪j���N���b�����d*�{�\�j��NQ6�����C�Z�YՉ����L�����[B�قdi��e�k�7�!��/�[�s��Y����U�܏i獍���M�&���'�'ڦ���Nl'���� t�kꍥ�_3��g�nW�f�_ت������V�#�ӸD3�����������������o���ȧV� i`��a�8�;��V-��$5᪶�V�1�$`�j��N����[�P�;�^o+����ו�Ti�fb"�G�g�k�I���4ҘuO� n�GcVO��unm��O/�44�A�a`��Ͽ������X�Uu,<M%[bo4�a�i��>��WQx�{����|�X_�^��H�@Ի�Sɒ��c�y"�F�	F8�-��p&И����8*A&�r�&�D�]1u�<��J�Y-N�>�Jum�.3>��a�R��T�%On�x8&��U����h�oET���)}���:��Q��."Ë�_�I�� ��醠����$U[���䨉�2$pPˑX�W�/�4ء��L�&�ʶ�4�

|[e�]�u��p�**<������i�Y��i�Ȑ��P�V�P���x����VI��[��&����(�����e���÷� �b���\S-K}�MÐu#/J�/�
y���q+�:�	�>Wߠ�����MC	�C'x2����=�h6���_>�@����O��g"6�ɷ��.���P�/�*�%�"@�(n��;(/�y�r���?�X̟�j3�u�����s��o��l(�^+j����B��fV��(��wi�/�k��9�B����6�T�k�Y�p=~���
�q����(�����|i;C�Y5A-��a���e����1��॥���.�H��򅙈��#�s_��p!��qt����I9v>�1�$<5����������d��ϚӘ���te��|`v"���x��4�D���=��Y�Ȅ7��b�x6�«��(�J�</�R����2��7"j����3M�u��)v􃱤��ڌ=$�Gb�Ib@r���"��Ԃ P��`��b���-I;��f C>����Q_�̟����(K��l�@!�C�ʷ�§M)�<;y-�YƩԡ��z�Nr��Dϳa,�4ܜ'
�(����s;)t��5~�AG�Mkp�t�/��x�\$�����/!$�������(�����S�VJ�I^���>�i�h¡Х���^rV�r��A9"'�m l��d��gϳV�Y�[:�`ka]��֍M���aD�2��Ax�\e��Yz�{�9�G�?30�L6��'����t��o��j�I�n$ܖ}����S�S�KFSy7�Q�9�pQDK�����?Mr1���?�p�2 �ͯ�"�dҠ��i�|o����ɑL����ۭ�)X���k�Pb�h����݄Y�ҹ�b��|�`��F�F�>FN�W������3�ɻo����v���J���N�lGkD�os��t&�Ul�g�Օ�@K�3����B)��/��v.���346�V]�M�������#M͂��{��&*Eu�ngQ�\k@�s	�ϱ�E��%�t�^��q��o�O��n��NО�LvV�{�D�E���`��}�Fm�;.˽�uc �Bk(jq��;�V㐸��敖�y3���z�H�*(���^�I}1_ �x%.�,�t^ba9#���W���y/������QI��P11a�,E%b�&�V�)����I�L��l�jS6�x�Y%�$pL9������h��Z�\�I�a�HpsϤ'�4�oe<u���u��&-_�u��v���@�*�mȄO���&e�������/�a�c9T�&%�(�b��y>[̿�I=���5��&�g8�B�@�}{�Q�(��"Kf������y�fW��%��]d��30B�X�i�N��r1��bE^�s���NXK��9	L7Y���ɒnA#���^�}��C��WٞϺuY�kO��dO2�%�0.<���Q�� �e���}������Y�ں9T��6p�"i�vܷ����C�����M��=M�Q�-͟����K��Bt�!=�c#x��W��F�@�!7��6��3,��Y�"�����]��TB�������������D�ɏQ��E�ƾ#��%��/:}�� �:.��o7�gk4,�X��_F|���� Z���4�:,@a�Y��%����?*o��#p��d;e��C;����n� TZ�{F��w@C[�kӞwa��A����YW��"?F�� ��2�3^��$�%��gH,:�l� mO��W(<ȋ��ܮ����pG� ���*���י ��k��2�r����}���� ��.q���la�/i�U��YR��&�G~#q��h��+|b\�!��m�R��,2��'/#@���/G<�8֛\�6��k���%�y��g�0T3�\�>&*2$�ow6����gO���^�ַ[:�!��SL�6�mi���ܢҺcOA��v^�WC�֊�C��;��|�u�}�Y�ٞ���QF,l߯��b��l2�j��+͏x��Q��y��U�E�l���B��q��{�}��ƣ��s������A5�E;Y
�D�.'/�ΏEb38ʵru ?�I$�J��`�:cfM�KY���4Ӯ�W�j�R�L�"�H�Ez���
]�����=BN�kc�>;߉@}\�>�/5\o��7�o����x�>"S�ܦ�����#�\��e�Tt*�0�j�����|aL7�>"?����;�G�mb"���!]�e�>kMt�ӯ���ނ��G��d����0�&-r�=wb��~ ���O�����!��f?��%8������Q�p$�ܒAbt�w�l�N�uX�>T�W�~�I�wx��ҋ��m�aI|��3���X@��>���tY
�,y��-k�l�g���y>��*]���1�#Z�O�!+d��U��Ӑ�CZ���L�:�V�+���Bo��2������I��u������%��/�#��X���%GЪ{��T��4�:0������2����B^�3����<�Q0���t-��A�F�;�|uK�gHY��ȑi��U�^�bb*7�҄G��`1��y�\�bρ�F���W��Zg����ٚ����-�^"'��I�O��BD�l�\�I�s�5��k$���͵�
cI�<"�qW��=~�I%�r)c2������i���~�+�
>�~Nj�����Ov�ٵE�s��ԓ^�7&Oş뷘�Dy���vJXu9��Y!���ڋb�eU����;��S��p~����y�T�{,��)&�fL�Q�J҂���as:.���f{_�Zp���af�_�1��1H�o0Fp1�rAF��,�}v�]�����ֶ��3��d�`�'- ���&yw���͎o��`�5ğZi�8��%���֟p�j񶙛�	��&7'F�	�@8S	�� ���� _e�X��	54���"��t�Ӧ4�n���!c�w%aj�+����I�(�*t_{�W��qS	���f���y���G>F
�Ҝ�xp�f7-"
�XFʮ�p��4P��ɓ7�(YG�C�ν�2���R)Sy��ia"#������N��jBynr��&tr���]	f@����U�۰�BW�3��_��v�掦�US�,�e	M5�[DD;uf�����4zC��I�`�)�W��㍟�� �=�}�Ʈ����jH����4����0(o�h,�	�	�v���B2N+
��r:/�jR�4	�O:�=��W2$�:��b`��ť��9��E$��ֺ����~_�6�����2��!M`�(�w�MfMH�ݮ,��Orp�x�M�0�|�1nJ
�o	�S#o�w?���y�
����͐�!pD�y2M�ђ4м�zҾ;\�q
pHo�f�Z��ՙ~{a.I��Xt|/(w�X��9ˎ�,|��R�Qv�7F�}���������q�5iY��V����_#j���Q�����d#4�:�^��)li/�#���ɬ�i�y��(���ꄉ�z�!wH�\�SB�= �(W(�EE@g�y��@^t>���äps.�a%�D�S4�1�qwXaNd��Cʖ͖�E)���S����jcD{qJgU��&1&�6�{L���G/��*�:*��y��0T%��6��fI��fB�a�
�ݡ�rfMo@�e���駲Ѫ����[3 �L�dT�g���p�xkr��S�!�f���]oQ5����2�`m�W�#�}C���i�^oZ�;C�]��&si"�)Ra7����+jq�P���>_�;�)��\���1FۡS��^�|C�k�(И�Sn�j��U\	���q�1�*���H�K�lf+h��÷���	���h+���;�PG^]s3}�3L�*����t��{�H�����Q��W��Q��A`����X������?��l���i��e����R�
�֕x�o�@�M5$����H�����f�o��\��F���e����}�3�~�f9'P�$Y�Q�Y1[�x/-�ޏ4B*k2�e���+�^��p�����s�Xİ#D Z���"�-߆�*�"�l��ghxf���P�C3�'�IjG��9�֯��P�&�����z&O�3��kΓG�"9���ύ�P�)�#f�XX��`�N��~� E��̫�<f�?�#R	���'rm�~}��L����U $}��1�	�$�2��tY�&�7(,9r�l��q�Y�P*�=4<� JH>�o��}���(��Ț`���n�jQ��UJ�ɱ;�]� �ިW8�zi����L;I�a�˲5A�u+eV78��2�\$�l�{8�ĚL�+�_b(�k�(Ա�00�>M��ȃ�#�����WҠ[��G҇ן[�\lJ���=Xl���^��yT���U0�G�9�%�D@@�zu0y�aJ�|�i���
��d�i�a��_�W�vT�x��%�X��wz��!�]'����<ٙ�,�զ� *l��'K`QF�S��~4�z��H�"���n�Z��}D4�]Ƀ������*M�5%�>:d�ޒ�y��q֖ϟ��G;?�63�[�k��洯��KW͓b}Z���tD]������.�Ef��P�����1�r��m�-�Yg���X��I���6�R��<e$�dz���7�+�dQq�g��@?[Q����.��oBO�=B�LU_J�G��� ���! oȔ�T��Mq����d��|I'�FΘ�6�k��Е�i��G�+f�t����@_��/�͇����ݦۿ���A�r��n�~��Ȧ��!I��e�4�ÉPX�:<r�yeNed���R���f����V�ƾ{ű���rm����LuS��X��U>y����f��;ʃ.�r������+���A:b4��cFr3O�ڼ��b䄁������+�a��?j�E�OBJ��#�;��r���gͶ�h�WZ��2��m���(پ	��dR��t��4��/�a1�o{��b�&%[�&J��)@�{�Ń V͓�<�G��^>l�HlͨD��M��!Ҷ����x�1ڟc6�'Lh���F}��[|6z&KL"� �7.�T	}F�&���5��W�8C���U�^���pb�mކ�s�i-V�����'g.��z9$��[3x�q!,���p��H��~I����ne����n���迥+Sv�4/�Θ�Fa�m�{��w�~�j�Luv�lɁz�z��8V�H�<�*6��#c�2��q}�����X�B�Ry(����F*�� Ǫ��s�V��2�ʺH��I���b]��w��r��F�T�c����F�ă�g����z�q��L�F"Rr��u��c���m�Ffɤ�C�ZD�����/���3��z<(]Un�c'ǖ��_��&�J�Lα���?d]4Rc�p=]����ι�������zt��1��9�(����}td�Ik��
�˖*s�(��F67<:�+�@�f��8p�o����K^̿+�aoT�k��bS/O��/�wئ�S?z�z���/�
�tyxc�2��O+9������iV$�|F���"�{�6�b%�Tw�)#�տK/;��ۡw�2��A��|ʵ�����.���b��T%C��f	8;��/q9��j�xH��΅ĕl��a>�[A�︀m��Q�U�K���A��,�g�܈�Gâx� lg;lA|D`���ө�=�]��o_�1��*� ����8+x���o1wI�K�(����k����m����_����ͣ�#��u��Giu�EYp�v����Uy!Z��1b�]I`��p-�(�6��O�����e̠���zW�D�ֱQJ�~݃٭�k��>� �UJT�u̥m��	ϓF���j��(�JPdU��[2���Mfy��G�.�!�@y�	~1᠃� ���,����K��~c����.mk��%���v�ٳ��:II
q�)�7(s���GAY@��ӄ�l5�m-�PT���k�׼�^<k�*�}�Oȫ�9۩�bEo�&�pa���np� � �W�����D�^jq�J#�5��n��5�iR-i�Y��{��4_���֫��E���叻M9��t��8��i��
����N����ݛ%��v�l��D&
��˦ΛV��`��X�u��q���A��4ͅ: ~(�˸���0��7L�1���}��]z��0^i/��X�׋d|y�|b�4���xT�>Z��� &{�;����W�
�w�yI�D	O���ECY���ܒo�o��ȶ�˨�t"#�spe�B%�tQ��#�9^JN��blv^�T
6s���{�r�aR�i���8+-��N�S*��w`�g��ǡ�ݛ����=�e؜j)mPީӻ�2��m�fA��jM*�Q"��Xaj�(E�8��r�w�XJZP�j0��#�mM	�z��i&�T.W�R�B�RB�����G���>L�(�^z!��N5Qzu���kw�X�iGL����>��'�ȟFжK�4��`jߏ����Sh�ry���'��Sw=�ы�Iy�a��!�B��߸���n���}ߌ%%K����T:BgܫL$��#��^��U��<����K�� ����z�e���!�=]����Y��D��*l�6���n�{Ͳ�
�2�O��l~6Whh�a�x,�������<��$b�3�0)�'���-��!�b�mw��#[V��h�o�Z�}���nG��V3��!��L�o��qdg�em�C�GXi���[����>�ҡhA���/�`�&�$��,v��ʕ�Z9�|��-���E���+����<�Ӫק¶>U1ݭ�W�6N癦nu��w���֤K��N��*XmI/�'�dj�� �eH$��/����%phi~��G Qu��2yz����P��)�UʳY/{�����ؚ�ͷ��$ǔ�[ e��>��r��.�6"*gs,V4��r��Z��a@H�P���}���S��{�nC�~Q�F���v&���X �~ɵ�ٕ���G�MP���H���G�"�U1%�t5�92��hE�㚈��3R�J��+-�����̒�x=�I��g?)��#)�uގQ����Q.Y'l������5��.���@�b1z:�(z�MG䄴o�#�ͦ���i|ty��TT��$��jL�6�,�[�[�"^��Z����?��6CN��Ә�{���vQ��}@�#)a�tAn�I�s��*�Z��
��N���-�	�&R
:޽9Z����&�UPnt�[օ|�����I����y���Ȏ�栚��F�n���b����,���T&��nS�7�*22�� ��^��~�ӈ �[Y.�ǳӦ����3��D��N���Α|��&d.�\���6*���qZKl�v�����ze�
t�A	����#� ��\��w7�]�hg�H�2� �.��7-��#��A�&s1d'l��QL�(6l��E�@]�s��U��g�����"��{h�+a4���G� N�el
����<��w��! d��ߙ����$4ׯu/\�5P�`Ho?���*CR��HI�a����D{i�)���T7�)>�����3���A�|?-R_��; �h K@����0�t*+�S]e�\����:��:o4�e�7NT�^�69H��$���r����DC�ʄ��<���f� -��`�����?k'35�i��j�@NP-���̘^?~@��2�|��!�c6��f{�YW�k��e�\�:>	�:��i" ���(���a��} S۩��a%$���4�Sb�=�e=i�y�e�����h#RqbM�=�S�hޜ�a3DvS׉\�
F�?h������_'�h��Y��ZV�|·O%�cK�����ku;;L��6àZY9"hZ�N�]壚�3�J鬞���!�-Y�Θۉ�o���OE�ΐ�K���&�J�y��$kG�g�7`l!�c���P�slk��D���}ˏ]t��l�X��G=��:���~�}���N�V<=l�-�&Z��xF��N2S�m�T�K�=4�UU(w譱'^�� �xvqS# �����^� z,�Y�Ŀ0q,����w���q�V	��r�7|��_�-5�ɧ��D��=!i���G>�C ����`�0sd�45�_����?5�y���N�ЙrK-�v~� 0�5a�O�֓)�
����ӎX�[B��;��6ɵ�������)(�I���ZMS���a���'���%��s��깰b�9��j iSzX�0q���1޹CN���#��23J�B��&D4N��Y{�wem<�Ϛ~^���\���Q̒b ϒh�����@mt般��{�|%�����o.5k޺�1y��#�/����Z�>%T��=�0޽����k�ȈZ6,��@��Q|��+��S6�D���x*��o�NT��ƹ����by_�̓5EO�w�"���C�GE��xQFJ���C�.������	������CnB�goh�6��P�m�n}1�6B+�ɼh��*Rl~��H�	y��*�T�I��v�,~��E;�%ͧr'Z'c�M(o���3�l�оUݣG�5�NmQ`P�L���:�8���ۂ͓��R�+;S�, ��W{�ղ�͸���1I�I�|�5���i����f�t����qޚ"��S��(�=k� 7f��(���.�@l�����	GDl�N�������3c���'q-`��U�Jo��Y�8�n�j�\d˜TD���ܻ����p�Ȫ�r��s8"	`"��cAn���~UU<f�������6&�����+O��D0|H`��#��I�Q)��WFG㝂R'�AS/g`��Za��������h,D{Xט�G'�R ~����k<���|1�mm�EKp�~ӫ#��_�Q@�O�q�;�ƵBq��TRG�w�3A�w�6#&_v���0�|2��G5R���u%�"������	�v���м��Da�K-�B,��|�����bYX�uOs�09�Ԁ&��;�o�&�R�H�|5��a�~2�{>x��Kj����Qz����������NO�ܾ&����Ώkz��� ��h��R��@X��s$G~��i�x���)�!%}��B�b�HW����8h��,�M���K"j��������Nl崞1]�H��dN�)7:˥:��gg������WTd��
�G�$� ���'6:H�S�4�_!��� ��v��Ë1�+]V�z>�m�����Im�vX��k��/Yk.a%��,�Q���Q���� h���GlM̵���vNf:�,��9l�D��D��M� �xt�o�Tk���qn$m���/H,0����1�/b��ι�ڨ7�6� e&ywѬ`z�i�z=��@��D�̺�r���MKވO�}�����tל����o�Z	�4U��O��Z��7�oI�G�ۈ��E���)˦8>��<�Mx��IY�!���Tc&K��!��q����Ek3��|��<z���O��[,(�	�8n�^~p�6���"������)�̋{�!�f�  ��>N�E��Jj9�2V���ɖ�,|��di,L�"LL�ow����U
��u�1�ػdO�������g�/��� iƍ���[{.���M/]~9?�Q�DI���p�� �$�^챬��fE�/�5��Y�����&����.ʔ��?K�?GpT���u��ۼ���gҺ@����[�g����;��3�'>�.�G�$�?nf�QF��ˢv���l�w\$"G0�V��jt�e����b�O6`�;�cU!$�ؔ��G�<�c쇽��(O��ҎƬp��;�=�yء���A�f�Z�j����<���N����8�j^y� ��UȻ��`Pf�`/Os��~��������by��Nh�� �7J�:�
���?\�!Sm��6��Ru�p��\V����3��-B;�l$E�g�g��Ձ�nF!��ۖ��yZ��r5fC��Ã:GTf�����i�?4M����;��lb-�i<��m��G�[�5�G�H
��s�l4�m�)��v��ۂ��"_�-q��q�a���h��@+6[V�'����Z�p?h��dN8�z`�`�WU䌓����_���ܼ�aڲ� X�/k���U`E�|�>�D5�~Q�'F�뭺k�q����2��t�Lֲ��1��o[�7�K+�8]%�k�A�&Z��ڍ�����ҵE�,�O�}��hKSzTo���P��
�^�ҾX��%��!H��I�.,���wڟP���J"�F���ڭ;�Y�T���a[T�}V?F��B)�l�z����igD�[�Q~m����c�4-�ފP#�3]�z�n4]S�˂��h���o�B������]�[8>�S2Fs�R^�Yb��k ~���`�iݕ�G��k<��ua�γ�����z��B��a뇤lũ�4��ׂ�/F�u7Ɨa��g�EaD�:�u��(#<h I�����Wej��?,R���XE�^�]�U*^LYF�٪�;Iȧ�m ��v��aj5?���iL�A����Y���׺=}l%y_���I��$0I��|�Ø����� u>^kDJ�-�1�rxp�+��r	AZ9>�y�D���GU���Q��^�r\X>k]����꼼�����L�MB���)'�"r�l"�U�\���2�4Yע�7m����H�@-Q��f��{pa)%�ϫũ*+˖�eE(G��L��� j��P9��Z��2��cb��y0qC�A>�n�D�qҞ<����y��/݋U���C}ʃ���	k��ѪZXz���Oc�L�����	��4�OT��EpRsY�=�R��J�[�RgՔ�Ϥ��h�(b]j��eB�R����rg��V��H�Q�R����DkY�v�����$}Y{a�jz n�������̶�$�/���wQ��Ȋ�-ꈦ1�����h�*F�A˓�3�!2��GO���X�F�Z�r���\9�,I��ȟ�"�9����6 F(�x3X�zK�BBnߠ�p0T.z�e2�� R�C�)�{���Y'D����bOjʹ�q���ڱ�.Ͽm��e�{��.���E*z��,��H9�v�0�o8�n�J���c$�Ϭx/&����J��[FhIbG��E&�sM<�olcz	y鴃�T�u7:���x4�z:��:Uo�\}x�F%�0f�b�jz@���:��'�jL��Bs�{�FT���aKoo���H�nt=�.�yt)��Q
���Y��C�=SM�̆'�v��7wك
^�t]��̦��3q��>�F�x5I��.ot
ݯ��b�rH�K�#Ң;��ȅm���6�t��K-��=U���<�D���=��'�łϋ�H���I��LE9ft��P��-����۽m?E�����KһS���}�a@�H����ѐߋ+Ϲ]����=�yB`(n~T���d�#_��p�j���r���F�P�Y��Z�����c/mAui:�������ԙX�,!��Z������-k���q^��fP�����`wޫ�/J��K�1I<x|����x����6��d3����I[�{�W�d>�ݕ�����ƦM�%F�] �?�-�&�oݢ�${d�e
�ݦ�c�LAH��/�%�c&H{A�R�&�'�U�'�[g^�M��q-�yX�}Vj��pc��2�z��OC�&�r`u�ɂ�|�/ 22BOV��7�'��~ZC�/Q��R���sZ�g+2�]�YP��N�����T���E���UA�
�>.�r%v��X�����P�pO��;5���֘�����AJ�zA4���t���ӺUMP��^,#��ӻ0�Lʸ�{�L�Z(���I�Vk_����țM�ჲ��Q�EIb?
 ��������)�V44��������+�Y[UD-��\�ܮ��̂ݫ�����bYP)8usk��5��І�5��[e��q��@��%{BFۆ����h���۰&�%E��7��%�|�z�m\���k�\�`�����X�/�o�O�eV#I�$�c]��k�a���'	��M�O��DF9��A~� ���,Z�w' ٿ�V��nd�3q�/ZS�6h�s�~Zs�����k��/���}�YZc���C��W��Ȅ��(�7N3�0c��'t�þ/WN���S}Q��6P�,���؈��"y�Iu:�fݸ�n���xa����!��~2�b��� 8�c�s{擊hr����9J���漣�4D��u@\̓rMj���(���vU�ʺgL����T��8�%����\𻋾f�&r?Dxc����n�@�$̏>��k&J�|�?D5�[��d����.�ɐG���X��J7����l���i�J�nk�L�3���f�;S�oc�廙�n��߸�G+I��#����iڴ�tDw��gN�����3�W!�*�j���\�'�@|WO��:���T|�,�N]��g�_R�@�1ǌ�������.�28��d`zc]�q��\��o1��E��n{��t�����"����Bs��?���ِ�
2j>Ց����+��fG�t�L�JcIfi{�~�3�Q�-�`�(�>Tnul��7S�Rù��t�����Ip�����LT��\�?�����9>�d�e�Y_+��E�Z�
�;byN"���߁֐ �.#�>֠#���/�;�!_� tH����k %�l��,3��eO�K��z#�v�'��ț�&���<Ë{�A����AZ��T���.��iȔ_:(�QQ�Ĥr�5���Vy2��#i�Fhve�ɽ�׍fgh	�R� �~]\>�_3n�ZЗ��ʆF���"����0�TҢ��bT��?F�V����������i��CZ|�w��4���sP���7���*	
��Pn_cA��y�J����Sm'#�p�k�1�~�I�t��TY��Uk�L����<a�W�w<Gz[D8�;P�.�n���c��G�(e�.�������I�G{6�%A�, ���?Z�4�z�GA+����������Bӆ�@t=r��ņ��K�F%�|]�Աc,����,t.��>�0�8y?_m��d�e)n��}+ ^9��v���ڲ�[��ű�+Ӿ湗˛����u�Ջ��y�1l����)q�� ɳ���������e��E�eV�]̞Qa�'�/4��=��PuܯA���MD��H;k �?�hQ�nha�3�
�3Ğ��u/�W�(�
�1X���<�����\C;@#�u޹#��-� ��2Y�ݥ�%��
dlZ�K��'�B���I��Rޏ��%��H�&�����k������Ȼ*�2輢^(L\���Ȅ4h�Z`����Wҙ�qO~����&
p�-��j���]��h{���$C�󛜚���*��-�y�t�?3�ʟ�[�F�(p��z���d�@E
�D�fCab���>�F���ɐ�V��'8)�c���뇧�sӉ�U���B���P�fL�Q�N�r�O�C�Y���P�\Pf��،��Q#��01���hhw.��qSL��fK̿��|6y���S�5��C���;�IK펮[�)gY���a<R�������p�Dx�1m��o����`p�Zz��$3�.����^�2^j1ߤ?�ֆ7LBc$_�6�J�g�6���fH=I���n6Q�Ǩ�z�mzo��-�ė�)���,�f�FszI*����&z��{�
F�c�mǛSA(U�9h�e�֛l0�M����>�8A.�?������]��{q��5��� �Pp��Y¹�zi/������`������&`2-Q=�(�6�+O����>���D�86ky�\�w��HlԬc7(�����C���!X�:B�p����|Q{�t <v�W.���[j���37Y��E�).�����qb��O؛�<1��N3����[淸�F֕"�5:V ?�K�ҹ4%s�F�%z�������PyX畫<"Lb!&��Gw�4��ہ���ZN���rt�&��ؾ8�.xu��8��	P�gS��J�_x�+���3?� ���yL;�*���ʇ���g�a���E2�.G__�8�����0B�m�gg���/�Q��g3��"eb�Kn���o��q�F�@�h�)��7���A�����1����ϴ~Xu��Z�y1��xS��Y�����-���j�*caNS�)���7��o�<���Q�J�x���������~��8P^��$}4����,:{�����	l����� H�t���o,nxwN�"�TL,P�o���ۧ��j@�C�J�G�F!�h�nXԪ)��3;t��đ����)�bGn��Io���%0=��Qi�k~�t`*������Z�Q���w	�ss��[u�� �����F?^<Aγ,��5�l�R�ts�e��A�@7$x�����P�������&W�W"�86��c�r��j�4Z:<1�-k��U-M�̌?ӯ��,.G���� �d����V�`�o�q��:Ǌ[I����ט�{�{��7�G[��ސ��嗾�8�<�ЇK@�!/[�4Xq�?��\>Y�.��p��p rsRp���6�A�?9j�����C�"����xfx ������a�WOƵ�
	�������B���χ�78�о�u�F�B��Ӌ��b�?|�V�9�	:{����^�Ϻ$۪畏>�8�؟��%����������d�����;�`=o�+TJA�B�K �߯K�3�0���8=�u
Ϧt Ce~M�;��J�؊�ڦ��)�.dp� 
8�j8k����̧��Cd�r�S�R�����&���8�/��NnWoog�e^�>�83�wm9�l�c�J�����G��Y�����8$M��˔x���֘]�
��te��M0�$#�o�f�u����׭�]����R+�%�a��>�`]*� :�mY��n�>�p'
5�Vf�c��GW8�+ݺy>-۽�,�ރL����W-ےJ�O��RLCF�j9���HvK����T�49o�� t� Q��_�m��աbT5�r���G��Gv� J8/)�Ⱦ���xL���LM<7m��Dl}�dZ���y�!��H��HK%���=���x�l9��1m����%�^I⥠��ѭ��I������o`�<�0ė.6~��,�m�df�}�f�L',7Jg̦^�6F���ҽ��>���Tq��gf3�Ѵ��j��íK��A��'`
���(^��dr1�3��k�Tj��X���g�/�l�Z�@�S�G��"��S	�����}�ߑX�E�ݼ�ˁ�������
��XZ�w}��I�$�1����x�1�mԁ�Q1����%.��u�#	�]�'bO�Q'gn��y!�}�J�a�l��}/���G�љ-D#���k�^�Qנ���`����qs>9�ރ�v[�a3�"���������S�sJ���^|�Wn��~�.�$���#t�0^�� v-��Qd�u�pz.<�X"�N��=i�&�����[�Kc�T

���k�|~۴V�3'�K����*
U����KH�`�<]�}y���d��e�_K?.��s
�V�����t�I�؈i��CUv�z�ćvJƽ�¡�g�|Ycb�Pm�����煩�/�9�mx$ߺ��Aڮs4X�STR��R~ �Qp��R#�:������ =3�o9�ɛ�OՁ�7>j[���'�P��}���Iˀ�ݷ�"�D�
���nYz�Υ�R՝Ķ��_0�<g�U�Ӵ�1�P^ |�?!d�����4#+�}�aˤaֳB��B^�q�q�Z�r{���Q���^�)�*�*5C�i����9��`��]��s�eF�������4��u�ׯ�]}��J����(��I/w~_n�]U�p�8�͆��p<���f�!�Q�+`��I�~J���B��0�:��i�׶����
�0@5sfv*�z�"rw�ru���P��=Z��\��wڋNrB��{��A��Ԝ"aԭ��@�Xq�S+PΡ�N�Y��{�.N�U!M\�] �5��M��lAi9�Ϛkt�(��/y��Z��~z��J�x�^G�6��#=7Rs��`�l0e���1���W�MP!m0@r�s`��1/ו7�0Hc6|Wj���L0b;�>3����jÅb�����cSD<�q".#5�����}֭V
#��4�I��*���s8]��#l��_�8����-��]C�U�bl��w�����NH�qe)����͎>�]A�M��9������E̝������Q��<��<~t��"POr�d���X>�
/�8uvr�T�J���"�O�n3�{�ȕw�h�aHq�g��WT`3能2���&0���5-������)��:F�֋й�SS�y�#��_��cy<�~_]�5(�qh�$�t�>��1��rX���s���~��Kȁ�i�	�Q����&4�a�?C�>.�c�����!�*��S�:���
�"��\�2cmqqy�+�P�Xj����������n�p&L{��?0}tN�����۱��Ɗ��Ƞ���2�;1� Ͽ�d|�\������k�W���r�]$�S	2���|ݭ|hl<IȨ�P���v.ѐR�=�/�t'޿7)�{\] %Er��:�u�Th_�h@@���9�/�1;��XC�����a��y�l��$n@�^��J�i��T���nYJc7�1��!v����m�zfb��^�T�cQ.�r�� ��i�@��<S6L�Z�F���G��j����g)kOM}=_S*���"��Z�G�s��K�c��P�5�����d^r�#
��2���)�邪�0��اu���CDx5ƉS�	��:��>DE�!9ʢ�i�N���t�Λ��ZR�J������3�W�97&J9����Y&���qۏ_�a0���)�����@0�uy\?V}<˭'[4��.�̡�	�߶"��n��Bu�lc��a
<�E���D�a[�;,$*���t���������{z��6�W'H'"	�'���DE5ۄ)D��}��j�����b�U ��� �7�RÀ42�;���mB�b�I2|#dx\^��>\JPu$�����8�V�W�\#�_%�h����Ӻ��C�>^�x� ���ux���>%�e�(�,ٸ�>:&ʷA�� H��%�˫���}��e�a�j+�8���g��ԗB�	5�2�86F�u,����@�wUgz=���wB�F��7�M�����z�p b�v&�!�_��i-���_����|y�Hu�ފ��r.�%�@l����y	�)b�6�,�BN2M���g��^�E�e����̨22Hp���&ʍ���c?V�H�.3y�77�-7��������U�$�FcbXJ�VS ���&>�o�Rk��埽����i8��� k�vz}v kۻ�	�w){{|�M�
�T�9���b
+3K�ի�����W�d�W�(YpfPR��������Nؔ�x�P�g�_�R6�>��"=e�	)껋r���5>u�C��:�.)h˕�D:Խm�W+����0@X�䚙�l����Y���%@�F/L_�랃ڬ�2:|&_�]U��8A�eZ�y���q�ֽ�� �����I� �O�/���Ol��ߪ �kr�5�ܑ��6������X�%�dN݈\��o��`�ک��[e�*��Q
�MPٌ�{t�[:MN�լǃT���WAk�'|�xs����T�z�}��5?�"�XV��?w�'� �|���$�$$�\GR�<�M����Mv��K��%�XމZ�V0�#=���v���VM#�>�[��O���S:�����8�z��0^�XH2�f_t���B�+^-����N��WO���)`�u,���1�i3���
�h�J�+�Kʋ�p-��"#�S�� ��2��!n��N��n�@M�`
����q����q|�2(�ē���Ls4O}�?G���F��H��cҀL�i�NuZ/���@)��X�S��ϔXd-�y�ǻ�:��#)u|P����cz�#�.��6�&h����g��2�-��6������|�=Q�g����%]xѳn
D��K�@�Lm�Ku����7�m�ȟ�Jʜc �o�'�{B�T�o�H���{�w���4kgy[���͏�}a���{�^
�=���A��(y�Z�_������/W�~/� n_�8�N�����´���k�����G��B�����P�/O�� N���w�黶.��V�_����07�յ�n���_[a$��7kaM���:��]U��<�U����+0<��D��m��x��k��V�J�&Igj[BKvb�%HP��R���T~�|9�z���7n�&��k���qsj�D���]���F��&ExFFz0��ff֏���w�g�#��`l�᳊H��������!�,���@�{�z-�P�`>0����w4�6څ�3Q!�3c��.�)�E�w?�B�D�fUΜ���z�^+/iem��@J�3���2��e�qA�2�P�n�=bnp�Ģ��@��vF�s��#�#�f۫ꌉY���.�[y����ba؏?s;���7t����L��vՐ�9�UEYZ��玊-4Cöjb����$����2 Re!�QoVAq���,?ڠ��͛����l�G"r��u}?m�#���V�D�[�+�Z�k�� �l�����)����^�rRW5r$�O{K:߳F��kLm�w!�,�D=���s�1.�BT&�=�e�/�|9�֗v��D�L�f��ex��4���@�F2[ �h�A��)�E,��-,Iû��8���\_���\�^U�d"�0S�&���7�k�C�� |k�M� �<�����b���!��L����k���a�M��j���L] �^�7 �Mh���B�[b�4x�UfVT�6#ɏc�sJ΄����Ɯ�~������i3��: ��c����X]�����[ �k��\Q kX	�"�/2�x�g�X�l����[F��Ԃ�`V�k��
�;�����=ӈ�e�+мJ��P
������u5ɐ�o�}E=��f1�e��%�O�.�vS)�I�8���w����!�o@磯��>��v�püu�7pd}��1x�m���{=+��$K�E�Ѵp�8q��yUj��坢�QEk���a�ʤE�������k���:'�G��� �S�o�Yh��_.� ,���y8�0�ޣ�����m.�����[�;M�7{�"�Iz��
�'E&�I�������pV�� bmc�G�,���gI�7���݆��(��cl��(��q����c��tZ�	�a����I�6^����d�X�p�Gl�>�|��O��H�<�3����y��~�ub�Um�U��߷�oh)�:
I���6�[�Ş<�wǴ���>����)ܭ�I�ħ0�%'&	e[T[�>�9$��ݭNյ�3�[�)E�e*���������o������V��6\��X�I�|��=RO}W U��W˪U�(�c�!��zVE}1���[��癝_��Й��2�
@o�����x;�o��s_T�i9�ɺrT��[K73\D eM��@⸣^���#&afUGmJ��l�98'4�W*�^���wG�9,񱅎.CK�Ƴ�U�Ҁ�&XtG�U��*���i���j`�=���Έm��"Qa�7e@ n��Zft/a�P��FWa�x�#��{pG6(���C��>A���D��{�PG�Al��˴LM��ð?�����f�s�ں,�
��3%��yyU��p|���t\��3������n�h����בͫw[���0��n��`#f�,.���0�5��h�g��K�^�+_n��>H��@h?f�5�U>�������H�x��wD�Tl�U䮠�˱d��Q?��C@Q��*�$&EOf�`����sq��]��BK�k����J/�)��b�U�/6�Ztӕ�K��}�qhĺ^��؏�N�<��ē"�"1:��&�]��ZO�Osn�HҾk�Se���9�8��N�v"BXjT	�THS$c-��� ����-���튝�A�C���Q�I�z�b#N���:�ˌ��{&rм�Ӭ_"ݳ٭�7Ä�i������x�$G�I�]��2Xe��S�� Q�gG�|8�լ�ല8��S<_UPhAΥE�,�b�H5Wa�F�Yie�Э~�l� :�<d0��C��`[��f9|?�.�,�k�$���¸}O�%�aCe�Fd���G����߁?�޺��� ^�3�;�4�ux	�ct�Rf�C���I����z�o<޵�GVݕ�u�O�p��ɬz��p�6��U2�!A�5^"����c$dk%������g䈠x$��]2lÏ�E9g�"GJ]o�~�.-e�&[����� ��޻��F��¹��q�=6��vϯa$�o� se�v���ߑ$мլ���^/�7��PC�r8�]^��w#L:�~j�9�7�g�*�qMd�g��"9T��*���?KD�1֮�g̛�3����`��'�R��S���>Jz&�D��&q�&�۔G�5�"V�ٖ��e�u��m��/JظW��ʹ~	<=%����#��sS�S�º��j��2�Q�f%ѓ�x�+⯬�=,hO�sH�'�JR?;���K���r��O��}Ч*�,�4�Ĥ;�,p؋�JwL�����F���;�3����S��1Ȑ��`�w3]ʣ��ʽ�� �㩕q��]v�S���.k����@�@�ZƆ�������6�Zj6�ٜt����r�p��Y���p[��PJ�V�#Y#W+q��7ǥ��@��%�kۙ�7�D=���fw�N���u� �
x��Lq(���K�bV�jn�`PP>^���e5~C�Q*�^�đd���
8�՛�+�}�l�e>��I暃>�])�Gmt+��|O�U�s�M�ۃ]�������55&�IZ��P-����f1/`�����W���vUO��pgڋ�7L~�p�"��:h�1j9"�v��sl��"f��V����I�C���33��Y|���
��LB���"�j���3�9ۚ9�@���ػǏ������
kV�P�?R8Naq��/���W�	3dM!'l�H!0>/���f
ϴ��ϳH����;o��ǬOy��Y%�K�����#�����Fa�E.T]�;��	�d�>wv˚�aH�S�+U�,ݢ	�h�~k����C�~z晖��6�B{,�Hp!��{�F!3q�̛��J�"aw�z:�L�.����ma>���(��ڻ�D��W�([D6+�gq����3z�/�͕}�"��c.���{�G����ۙ�e��O��p��d�툔؅~�w!4؇�8�D������ep��}��ᰗ|��I�#A����;�B��<�$�� R�iSu%�W�s���W��?�z"��1�K�$��P�FRyT�A4(D��e7K����b�ogr�=$a(Kd�&z�����B���#�#U��?RV�������[�o�`��S��_"~V�h�{Z����C�Bb`�|�y=�ɕ����7�L��Suߊ����X�|!��c�zn��̏�kY9t%�N'R5�G�#�}�	���Q���E�)�e��k���fJ�����v1+��i�J-0[��3����JYJ|L�����p4"찳\�C�(ۙ/.�{O���'v!�����̆c�3��s����Q;^,[����1�2x�~0)��U�S��M�	���q�Z�c���<�04�C�FU����{'P�~!�BۙI�)�X��2^����s��;����ҁ�-:�Z\A*�
���e��pU��H��L����F�?�zd����`���6��V!�b�WV����;E�yק�W�{^��,u�n�P���A�,��V�pF�6�a��3S�\�A���uô7�Ĩ-C��0�Q��dΜ	O?2w1ٚ�����{�(����L��Y m����Č/?��P�ML8��r����$���!s��'�қ��!���Q#����� J�%�xʑ���;"-�+�*�6�z���i�^P�=��E���2�WVgrG�0�UK�dG����0T?��eacH��4���T	��u�S�X3/퇰��~�'mՄ�����B�b껕�CE՝��Q��I�v0	��hA�4;���<�O���{fsU�'��P�B|������w��CQr�����(���\�'��-���u��F�q�w�J��,Ϊ;��bTH�5G=�}�vo�����~��Vh຋�IP�����㜍�Պ��4��:t��R������轶5���/t��B3���*N%��U���<����3�1T61ߘ��4?>�0��D*�'Ŏ�8o��ء��9e���yu^G«�W���v�*q`I�e�C's�I#Jy`-����?5<��v��E��)4�l��t)@^`���v�}��'Ry��C��]��A�/�X�;c�{�ks߻Pgf������P����*�w9q��;\�����n�V�f�5��gش�|B��3r����W��r�����g�~rR�l<��X��bӒ��N�^�l\s��A��B��º���C#��ۓ"��d�9����z�+]8�"'�MQ�A�dl��R˚��)�+�W��د�U�S/�<\KK!��ا4G{�x�Y��x�3s�Lj�X�\��	��m3�K`�-a���WFN:.1r�3��#�� ٓ�=P����6�bD�d�w�*�����(븃2qAAc�=�d]���=3��[Xj����?�oc�]ɇ��-@�)��7L�D��!�.�5V��PO(>��:�;��W���3��˅�Y��R�˛/B�5xni�}}�~#�aSU�
	�7��^��W�E�{��E͘���7F^��,�c�W|��_��VO�PC�q�=�^M2���[2.�n>l���4] ��W���md��;��z�N�9�mTw.T��f�U=�d!t�[ӓ2��+0�,���]�&T'�yi��p!p�ZyVaI�)�3�s����0�H����k���k;��ܹ]�%��Yhz�����r;��=���GM(��AE� ���_�=�ZIi�i�1�N��4��0�L-dR�ΚQ]Z
6t�%�8��0n剭��M��֭��F����/��&��G��ռ��#�2��"hJ�y�4Z�&-��$�#{�̠�M���?=68��ϋ���|?$H�up>E�)+�$�vP�ݣ�ï���q�;�MLË\�Y� �rTE�
Fmݶz�J�d��284��l'1*�9��3���3
�,�up�d�쌞�A��m�Y�m���o��W��&^��aiނ�#�|�5��x�P���cN�T>]����j�]�����1������:g�n<jh2A ]9���)/�"4f.�����^ $�t��'^�=�~�Z� �%QhT$F�h
�%NE%�l�]��]B�A��*N����8YNL�T.�v��թA���ҳ��%u�?��9�W�:Q�.+qn8��M%�Fce�DS7�)e���{���0�g���R�u���H�π(I�hn�vEM�4|���� g�f�	f��<ZoY�������߰½��ef�~�`��1+s>L�~�Z$jAP�\���v��B��v~�0���*Gy@�<e��������s�̃b��o�ιJ���nIХ4���M�ҷ���%�1M��c%=��od�(�G2��;��mi��]��xhΰ���0�ͯ�$�A�8(_ѳ�Mu�:����>z�/)AÛ�3w���}�[��|E��x' %��؊?a.��u��:&��f��_H��X��(���p�9�Y�L|0�;�4=y.�3ۅD�u/lS�"U�r
�wh�m�{C��у�6�Nu^ڜ�yG�[��8E%a}I T�c��d�\X1L����h����R�_�>��:�M��Uf{��#��c~�j6c]�8���l��Bd����_���a=�o��߶e���b��i�)�&����Q�����#��m?��f[x��%�t�(��*�}4���f����M,���zo�"zC��|s%�ղ�)���ߚ*��[	e�M���!�������������u:>�J\����K���*�|�z�v�6�[��3�E)>N�Gۻ�G�򶅩D1:᪁����f�4��˓U�ہP�*���vg:�xXw������O^����&�or���#���n)�S�yd�˜�0^�.`�\ �����_$VaSa���XS�aﱁ5�,z^�ש�a�B��ji���F���+��|
�!3;�7T���}� Wj��UDh{W�{���
���	�a�?���洐gHKPo��͍�MA���A�ScM����"�=N	<6��
��c����d�IS�i��bw��j�@ )�!y1�:z�%�8�ME���*�~a\�X���;=Pj����O�@��	K�=�WaL��i?Y��W8J_�0�����?d�<Ik���UҒ��{I��8�[Y<0q߹�C���m�:o��/��Ie:������Pn�cA��
a9 �=&�� '�/�i����'�U�{)��ũD5V�U��ү�EǪH��]��U��.���m|���xr�(8o�w5#}���j�>�)X��x>!���m�PfD�"��!ni׏�L��gL��n Qw��V�n���j������^�lL�mk�jmw`hSC��_r���b��d�A�d
5��2ؙ���pҞ�����N��{3����қ�L��Qw�>�_���&F���K�8��X��+wK�,VL��%e�B} trR�m"G;˳� �R�j{M�j-�2@���i�C��G��<p�J;�=pH{,�'�"�)���v���o/K�W<�ıX�{�������f!|��OK�&�����&��bb�+]	��d*��<��VP�9@��Y����WQ33��'й̗�?�~�cN��q�^��2�?f�ǽn$x%�����$��j�Ih~���c����I��[m�s9�A�*$:(FV��@�_cg'Ҿ�)�\.1k��Nϋ���]�6��or|y��H����=��>n��Yc��vۭ��� ��4���-�������S�e��u�?=�)H��ؼH�?�B̊��J4��9oWiIR!j�/ʓ�x�����b�"�l��w@HN*a�&�� A�܏����o�g��h��q�M.5��f� 	�@0ֻ�ҁ��L�y�1�fO��E6�@���el��c��0�v�Px��'�nW����TEŅP����.<��!l/wSL��IZ�.�˵���,q���>Y"L�6.�ԃ�p�'r�ҥ��7�h�3|
�1n;�M܂�kf�%&L8��_��>���fu�x�� ����[=cgn˻��E���ߍ�!���wT��YXft�3]���OV=0���C��G�<���mo9�#��p�oUi�M`e���I�U���:*��	�Q�2N��ı �`��$;a8UG�~����Ukp�y��S�k5�ر�{�G��n�T�3����g������`�R�Xn�j��|��@�<���S��2B�
"�v	�t��J�[sB�2%Cˡ9�(�8����5���������coy�Z�3Τ�� H&��7*�jzZ3� �_��$�r�{cr�EB|	6���e�����U[��e����z9X��9 m�$���J��I�Ǭ�BX�Z�΂];��D�K=#x�㰔�.����E]�P���Y��{�y���=�d���9q���+�� ''���.���S��9g����A,/�~�����Òuy��m3����;8u[���!hG�dA��́!�Mٹ�M���?���:�̡�S�a=z'mZ-@�f��c�0di㶆y`l�����Wo_ݪ�h��S���;�ad%�G@n3�>)��xv�#��=|�"U���u���� -�q_ong`��d)�bWEҥ��Nu�����ދ��0I�H���9��nz#|G��$2 �Ɨ��gzl��y�@JJ�v��c����$����xV�)��>؞�%6^B���&X���Xk>}�]��R"�l*Q{�N�6���Y�R�Юw�Y��^,��oĥ��:́��3c��=�sj�$T��w�1-c.M��!��Dd�z�h����)a�c��vq�y6hF�f�*��e���{f���@��4q{��à]7ٸ��)H�<�+wO��i0����&ܠJ�'�<;�rk+�́�U��wX�>ƾ*.�J�1kjBq���V�/�!��b�!;L��N���0�z"Gl��X�@i�;5*�$��(��^D�c	���q�K�qA�79ybwO���`�g�v�V�+���pDn�CxR�=G0�"�(S�N�����P�]l�դ�����:L���b�?o�Vr�I�E��v��G8$&h�,g  9�����g�Eن,-��S�E��������<���j�6���n�d42tYAˆ��mF�b/��A�\5Jݜ�t��\�b�+H�����<`%�4"�"�nD�Uw���]��(����30�-e�� `͔���D�|\]w�V�4 �c�s�[�p�p��2N���'3�m����|�l�RMA40��yvo� �%��|ƨ	V#
��"�d�>X��G�:��PKC��+��W���pwI�ub��*Gs�%A�!z����`�q_�1��QtI-�U����Q�Cm�J|�$[�
E�������T�:�I���h��4�=��}=�Z��f��#�Na����:5�\�{�oX]5&j@�����t�<��������N�d��d\!��Y��5,ި	$Pt"�^��w�9Q�t��H��R�J�&fs���;�_�E�6�� �7�}�������ց�}�1�2�1\�@�V���rS�~�dφ@?U@�-��v�ʆT�/W����tw	��	�u��i1�Yz���6H�L�	�i�	%3��ר���O���̶�@��ŷ<U�ȅ�;ҁ��H.D��'��_TW�I��k�d3���P "���N��>�baK�0�Z�a�K�)���ݑ> �(�o����?��9?P�q��m>E"�TQ]k򜴹ӎ�����'sE�V!��;.����>����jܩ�?ʼt��O��_Ǳ�z�fv*�1���Daƻ�"��hޯw WY���u� �-�3~����O�����f��&d:.����V�Va��<��S��_i���w�{E	qOxb�Ra�M����!��Nu�+8�
��P7���|�m=�
Z�d3ZM���z���:�?o1|�8��/�Z?7��L#	�Ε��ɬ�e�%�;�F��<ހ�00w��
4�i�N�x䫼��`�OXp�#E�>�#u�2�~���3��l*���n6}�Fف~,P��M+�dI<>8�Rx��*Y6P ⦤K1�>����'�mZ�ʡ�K�1w��m'$�?{=b�/_8R=��V��^��jH|�9h�����v�Qr�~�,}Ѣ5��oȂ{� �M��H��o�7������� VΙ��U��#Ʀ��oY9���$��g,+��`��5���s?����f�؛��}��w�����֠HԞ�=Eo��p�-|���ٔŪ�����`��mxI�X�UN��^�Ǎ�@J�5s-�
�y�dO��SE8���� /�~�<t�z��B�d�+Qɢ �\�6�x�D4pj�g��Q�h#�ɘ1(�г3�p2[���R���ϣ��;7�t'���T(��I�4b�\���fL��R!��!�\��Я%/���/�bT�$��;��+E9����-_�&Wǅ��-�� �,�s��  $\}�8gM?��/܋t�`�`r�=��@pu�*�M8�^��(N�6=��QER�e5��p��2)�w����x]gD!s�⵪�l����f���8����h��n�CKq�f �֮p��0��l�>VHPzq'̬X��n�?$6�=cC �[R:�Hb���nAT�&��.
�bYx��at���b��au���[�tH�p|�"�{Id�~�rK/D�P��Ӆ��4���j`홦��<����<~{�l�
�?˯�H��|���F�Uo�w�,�?$�������ݭ�o{�/ȸ���&�S9�{}!�m�+{�e�ꂣ�,�i�5��ll�ٙ<�E��m���k�zތ�HԽ,`9g�x8��m���vk(`p8w����=�A��r�����Kr�ɀene2��8�y�d�h<�B���kB�N<Y]���G�΂�a�S�^�υb�u���S�2L��g�h3���~=�-.x���saL��$���q�J*3�Cc�Ys�1���e����M+�Z��a��_[G�X��.�"��%���'�@}N ��'N��b��sF���+|�x5��v�'��J^�O1e". N���8�z����?����?������6�:�C��K$�~�����$�7���`B-Zz�ѵ�JeB I���C���Hf2:�B#VN�����ؼN�9O�\P,A���h�[e�2�L�ݗ��`���`c\.���PG00>QĠ�w��^����J;������h��dGaL4�Q}��cP���>E}ͧ�}�ή�����QCQa��@b��^��c�y,�i�q���M��b ]��y�`xx�v3曤��_���E�75�z���x\S��a�� РL�������,W)�/۱���w~��E�}�T~E�I�V3 Y�i����9��W�˴$�d����E��p2V'��T���*_KnU%9-�K�u��{z/7�B�9����`�t~�r(j�j��4�>.؁͠�_$���HhNt��_�EJ�@�i4I�ְ��'���`-����!���tP�&��Wą�v�k�TP��P�h���1���l&��守E=�)����~�#�Cr��H�b���U[��b��ݱ$֭�X����{u�lTҺz��8��"o�UO-����Z��D]����]����m3e��}�HHÈM�u�o¢����ɘ/f0g�j�/ua&/�yB}0@�����,}�NI��y"���B��zBjD�����{�u��@�M�)�Ɨ����_7�2�(3!�,y.L��r���~�Y�2�n�����zeb�|������R9����Fh�`I(�7����y�g�k��.���?=�R,�AQ
$�?n/�)���D
�#H^�N��i����(
��hQ�T�J��3E�'���y�������"5�ɵr��������o� �;�?H�z+v�k-��q@HѨ���W>4v+��~IZ;e�ܔ�/���j��VAϔ���pG�U���̫=�#9��H){�����!�[Q�.C�:sڔAT{��M�D���WJ��T���)�瞊�g�o��LG�O���4U��i��� �S���X�u�
�K�����S����q/Gn⃏�gz+��$�Ќ˷N��5Nh$����7(Ŀ��lL���j�<����B�S�#��I`��{d���!1y�}',f�չ�p��K�KO��s��庶�=� y��<�
SY-d ǅ ���MbU��$�ƶj��3�Ǹ��V��m�M�>����V��?�wU�pf�0t�%г��.�sw���I��b)oe=��Je�ܓ�`/��)�]jE%}�{�h�Iɑ>n��<i�З�R�9�R%a�M��C�j��͇:�e��N��|L��<�	�X���K���Hp���l7f3dp9K��v1
9m
�j�/6��`~�K�;^I�D��~R{��T��o�{����5�!��@�د,%�s�hѻ�c�Ata�~�sW*/��<GĄ�\����]_k�����,��8��/�|��� ��Ch�*�<��ڬP�g�?��aZ���x����@��Zԁ݊Y�LE����zP��R�^Pi㚓���e�ȎІw��NgF�2?h�Y�/e��C�Q��?/؝)k�ǩo>���s C\������%�j�Jp'�rf��;QqO��_{S���$!��M��ԉH�o�~C�~ ���V
)�o���>Il_�'���)?�v4��T^q	��� �2@����6=UsP�Ӑs"��e�@{Icak8 ���f�3����|Ț�v���U��0�S_�vxP
�������i���R%�'J��h����
Y��,��lfF}�=��+�aE8V����O��'���QE*q�?41ɾ��Q8��y$^�l��^:��f9/IЫ!?&o���z�A݅�}���=:Otȃy�Ԃª{sUVK q���F0b�kk����Ri.L4�!�T:��A�?��޹�*�L��D�z}�/�-l�
�S[&Őo��?4,1y��ʂr�
(:4-W&O�ɷ����Z�R�b)�ʀ��w�*gJ���4�

�Oic��йAhp�r�]ٍ�
�0'i�]��/A�.�$D�hVu�r��(!_<�U@�-+�O��0�sC	���c�����@��Ӳ0�5���j�����8����lMY�xX{�2RxL�Tu��:�0fPyם;���O�~��N[��S��a&��;dr7���<��йV���8��~?Ms��Y�,L�vޑKyLJ֋�C����2�`i�b5�袆*H�>8=�"�,v͞�}F��E�i��� ��7��i�.Ӝ�cZ�k����P#bf0k�V}]t��A<%�ڟ|����D��x���0�#�K��0O3�_J�hOr��?2�=��Y!hXȦ�ۯWt��h�b��HO�iv��=��~���&����f��������s@�>5ȯ���;�>T��zvv�?9���oY�7	�!��D?�R&a�8��o��B��7��aiݓ��}N56Y-�'(�xEdə���j6�#S�ݐ��4r��0I􁞮E���W+yQX��ö�B-lU��)i,�:_�g�|��a<ylx� �$$�y�����E�Ñ�9/ܚ9��Rǫ�h�������\�*⾒�[;��k%am׹3�(nz�Da���a@�luBU#�*BOE�u���1f��Ż�9�"��M�wm (��;Ygܤ2uz����gr|F��&M����+������NZ)*�'�3s#��~��$.�O�z��$��|���~�S%j-�YΠtV� �0��9�H~"�H8 ��2��!%�������O{�jn�h��F�Ss;�E�e/	bzP�{hn���.[�TK�t��_��q>t{M$���v4=��5��v��t��o]�[s�܃a���OUך�0��2�ML�'�F���C�o�@�$�;53�R�6噐�.*��Rj�위#��e�p����#�S~�Hs赗���@��ű]�_8��W%����dX?���nF���%(GjU��_q8@�+X�S��.�{����sEZ�����(Ѣ-��<V���0~�%k��g�ؒ��~�c`ȇG��Εʩ��G��6z���f�o}��n �,Õ^�+e��9���pW?9oaOL����F��])@���H��/ҳ��t@��+��JA�+�����c�������ȱ�#�n��z(9~��DZv'کX� �M}0�]���rϤ��
��9uMv/��;N��I�s_5���ٵGj�@�.TQ@#�����?N��G��s���Xo��ہEP.�oL!��f8���Ӏګ�, *%� �0 �lz6I��#��O_�H��#��-��`F;�!���1�9:θ�Ν�Zǡ��Ϻ�ii�/���o�ٽlyBk9�Ta�o�5�&�S� In��w���/irn��xD?���j(�	��	2XR�I������yl3��8����A�^GK��6��U@F�e�]�-hޱ�	�D���)Bβu���G�ƱO&��b�7�?fL�Ph����y2J��fx �u����E�,��%y�MHO.�J �T��e��|���J^���Iz�,v|�;~HN��C�>��ذ3���뫝X���U����f�	K��4�q8Kf�8��λ��R9�������
�蘉����H��_��қ�I73Q��h#ܵ���1j�Q���t1�_Ŵ�ca������D.����	�Z���+H��B�L���Z,͂��4r[;�&:�k�1*@�5EU�KF!�ğ�#Ú��J��h]���;�<a��Q�.�� (�+�O�-)�Y��;FJ��Y�'*�R��Z7�Gb�Յa�k�HC������"h�K��&K�;i�r�:�xn�s������=)�.C ���1��{H��F��Rc;�3�?GI�H�PZl�n�BP��=O������`�ܱ{�
KP��c0[aA�����rв��߷��M���48��pl��Bt,_/��Pt�^�uRbʱ/��;3K�Xj�?
�kڣٓ�C���t�ʑ-j��M��aܠ��GX9�����.�$z��e����M@�"�B�����g9o��/�'׋��\�T��ԅ�����a�<�����Ii��(�p�#�m��N����j�����!�@wV�PgTy)���a!nII���έo����Й��1��t�V��
�h��*�I�%�u5�z�U���������T���xm�ʽ�o
���7y��G�%��׊3al�#R �?I'ٗD?� ��WT��L��A���1�4��V	�6JrI,`E�����e!1\Q�63��?����:���o�9~Pa�],S�`����A��Ҋ���֢x�����
 ��g�R%�]�c=���B�����>8}��ϑ�ȣ�����K�s��5�)��á����n�����t�0u�Φ���_s�(j':�!}	�f�K���U�;F��2�p�AsCҿ�LU�7��G��y�C�G1�7�^rty���MY�:�=���3�^Tno���b/�RQ��Z/E�<�D�|7
^���T�l�/��.�}�\��`��V��1����)PU����{M��BG�4z8)�b?��`���6���K��]GH���L�G�|�Dۗ��4dO��Э�G�@���v.ሣUn���i��wt�=j|E�#�(���3/�	F�_ORq�e���2��[�1h�&���u�ɧ�>}-��7�qe��g����ܪf�=�����ao]�`*^!VM0������F��DM�$������	�R�%�sb[RI<��>��!��L�9���y�-ǌ^�+���>*�<Ze�HM�����J���ݏ��'&i�=S�]�9�g~�
%��©ZM�AKӪ�9ȥװJ����m��TJ?���&�(+_UvS;Ž͑����ɌoЛ��a9� ���fu��پYаXhk��R�j
J�V�b]o�X��|��LG�^]��s���T�&�{�h��A%Z��h��l����;[��7��z��K��!���P M�be�<�b��nPt�WM��$I��!I�Pcۥ���2�5��?T�Ɯ 5h�*����0:;�u�Hi9���ن�b"��*F2�	����i�+��g������!����O�@��E��م��>��ܜF����:�ۗR����n<�ab���{�����o`M�{��Χun��=�UD&���*�g��(�|���P�G-k��4$��|;���#5|"!P9h�-�-�}�"&C!3�>�Dh��wŀ-�d���	�i�[i>�x��(7_�E=y�z��˰%�<�ڦb&_'Ir�Az1n�%��T�s5l�N�4��(́��3�Z�9�(XPc�f�|`5�:?e@ �Pf�7�NO8}�&t�R���j�e:�u�0g�'�l���&T1��;°��#�
�����;�힁�,_�FƬ
��jd�l�������_~1Q_�����X�D�\�u�Cܞ�Gt��&p�{�+���݌��a�t�Hj�	;�~G�k&D#TU��H���	?�9_1�*�����2Β��u���q�K��"D��D�:drC0	��p����0�J�4� 9,���p��ܣKq]�Q�q-{O���pB��4�6�w�-�[Z.�� ��lU��R� �j�� l��9~��|j���t#tn:wRI��������x������tq��hmR�I����o?R���=�H0��|����ԩǢ�a�,@
"�����jP�Ztk�� �r���l��pu�
�$�%�1̶��89�p8����Pm��x�9�Ů��ic�P�^":)�m��ʃ1��"ٙq�A��6Rª���YO�y� >o
V�E$�ԃ5*�Kmu���f�0���z���qVu��1�S5�ֶ;�+��f�U���O���6�ҕ���p	~��Җ�n���w�����)ݥ�j6�n���,1*dn\ʻ�M�j�w[�Γ����[D�BP�J�YÆ��}���w�1Ts�%"�|-���g"]���9j[� ����a�%uZf+�2�17Kc��0'7�6�q�r��v�4�emx����o��0nX8'�M�f���>8�����V���E%��sNF��Q.
�GN�o����.���~�ɇ�		hKk���Jg:+�X�!�j:�B&tW�+��pd�~.�LO�@f�I#�u�"�G��2���p��1d��C"cr+�����W�$�u�t��q=��?���=Moz�?X�K{	P�����$�vd&i�;�o��A�e����2��p�dtk�u���h+l
�ߒy|�.�L<�Q�_���D�y\*�,������b�Q0���Is�.�:�d����
�o��O`������To��OB'�����6��GZ������s^妦�@��c4���mo��uX��=��L�-0܉?h�<���k��z���xt~n�Mt���K�c�v�v;aLV��s�ʘ錘@Er6�3�� ;��6�MƗ}�@k���}'��O�H��}����,I��8�P����-D��~�D+�z�ަ2�E�8��Pv�Z��nZ��S/��G�*�p̣�p�Q�^�A�=�����`?Ƨt�d��j+����5�G�gō��i1��+ވtJ�!������|*哂(<<�ڹ_1;�޸�u�kG��u�ܠ���M\]���A��[0N�9ƪ<Ѣ8�eKi������=�\�/�nhe��fPW|��L'!qyn�Rr?���n{(8k�>k�e�����J|��?fK8�y^�ԅ�N޲�(�&Ћ��/q�0a�3���<�]�;m��F�T?=E�#�����j�v+AQܜVRu>��2�����D�K�+��"p%���&���"ߍ�e�B�U�R �y8�Yy:Uotu�I�G�H��{���y�q<��N�n��qRW$���	l�Ђ��~S��f[:��G�:Z�D�i31}i��1`#bw�ajŎa�bD��[��δ�a`��I�^M�+hX{3R��G�\7ശ�m`7)m9u�GBg����]�N|���D�{�|ix\��Oo�*��Zue�m�o�+�*�{�l�y��� ����g�IU���}V ��Eg����>t��0o�ߥ���Em0{���DD��Y:A�Aa`<�95���B�c���ޘ�k���L,�\�	��5�3�
���#D�]1����f�kz��Id-��2r{8���£,;@�7"ԱOQH�'֛x�"����'[��:�׈�\TI�$D�]�r-��ȁ7]GT��U!��P�<oaA%����v�:����!�jXzn�y�����DFN�a�A��fh"S�;"8h#�5M�TL� 
\f����:��p��9�?�'�'E�hC��5��S@�M�48$��(���P�"�x�(���]Cb>��mI�5&6 �$V<nvx��Qq�=�ݕ������qe����>ǖXi�ith�����E�P매凩�&FL�&+��Ǫ�\Y����[Q�@�E5�Rz.���� ��\���J���������b�)`</�ކ�«�9 s"�o���ۜ��$3�21���15m�(E�sӂTAR��jǎ��t	;�Yt�ׯ��Fp|�iP%f���]�<���|�>�=����ې.G`��П�sS�C�����fP~��&h�FO�Q���N�� P�V.�saG��k6B^��ڜ��h�US����2D����r�A��l{G��	i\c����q��R�6}�����*�J5nt��n��x�
�~VjL�O9$So���b���Ӽ7E�U^�YCЮ'�a�$�����
��/����9G���Zk	 /�F3��jhIq���s�.����ｙ@�C�Y�f�LS�|�F�Rw��U*�Ч�����R�6cg{��4��@p+����#N���-���L�"��;6S$أ���'���@�8���/9��?Ǝ�'au��,�h䭴��&R��i�h*8��}�&��7Q��?�%��ٵS�(H��}Gm�ʚ+��qWIJ$�%�1��>扰⍰��Y+x��#����D� �=��[�E=B/E���YFy�DQ����>�1����p)��.�oi3]�dV\�3���-S�=u��'Ȃu��>Ϧ� `��
�i�bM*���q��n��@N<��w�3�zR2`���P 5�[��l�u�x���m�Nm�^�}�w��ɪ�e>���%�R�9��1��=�Vh9;߱O����A9�EE3s���$��+!@N��1���Ƀ�0�I>�^���P��͇��$ݬ�OX��ܒ��@ �[?�����ÿ1���V��]�t07�N�?��=��F]uY�7��Z�T@֊	��)z]���Ȋ��3����h_���=��X)97�<�q?�� {���%cGX_�^%Nw�6w|�,<��F���cI2auh-I?ߖ��ᒺH��dE���G���&2��9����#:e��Lj��JM*��#��m�hȊ��_.)�v!T�� gSG�� pYS����P�<�R�+� ʎ1T|p)q��7�ug�B8ȴ�í��gl�5�(��1k�81��9�ި!Z9O���v-u�T?I�
�����"� �u��Q��\D�S�ٌS�g����Y7��ZΝvޥ29��?���6���m���C�!J������/���"sVU�)��������k�<�Y^[`tP���2�+�Qc��k�?!�E�u���G������W)-���j�/��O��Bz����;�����xhz!}�_B�1?#{xky$�E�0 O=-��x��čq�4R�)5�/�=!-��Վ&�y���W�8MZ*�4
��,��'/j��/O��X0 jkB�����ȕ��'�-��	7��bjn���=�i��})���N�������j��"�2�젍i�ć�N����3kp����G�����Qb�1�8��o�$a�u�À������7��w��p&�>g�5�k��A���;U�Um�lyc����Ҥ���D&��_�RR�L}��.��\YӚ�3�	��{��k�<(&B�ϑ���ҝ`Yf�XE��2��I����_������
6��v4KgI3Y��RE�KX��^� \�P\3}����M�@;ٱSTp���� �
ٺ�"���K��z�JQ�U��O�G���_�۪����M���>a\��-\�.�x �s�P
UG�E�j��K��a�@���*�V:����*3��	GX��=i��U#x}( �T���,W�����@�|ϼ�Ѝe���K��[i��.GZ�USV9�
q����/`�fB~
����Ep���8��Yf��]�?;	����V�@l���H�o�\ݹt�7�W��`K�ҟ`Sf�i��ء�E������nbӌu��1��kͬ�\��g/�4���%!h����A��	&����:�
)����C>�+GǇ]�s;�`�΃^DlK_d�,t��+���i�����T�����HD�Y�����5�*�}�9*n����L!�)��"�c�~���և�/p�$:��k�7��Y�[�����.�hO ,j�H��t͊:���h��j�$OG(��.����oP�wb�紦�s%��-��A�a4��K��ﵴ&��!P�*�����Մ��'��J�s�0�G��n��_�Pj&x�!�G�����:-p���ԟ#�JTNj��\�! SuYY���?����FF�ނ�y PU�C� ��;���H7RO�uʯ/����n��X^$�g�+�b��xa����Ũ��38��Y�V���v"�i�=Etj�~15F2�z�!�9 ��RȲ7_!���C_$1%Z/W����}���xW/9�;Ji�<�����D�cM4۾����K���	�dM�٠6n��Q Ѣ�@�Ө�=��/��6�0�|�����7fŇ乭�:���/��
x�
��#~���/�ح��Y�6t�eKD'�q��"2���v0y�~QGۼ���}i����v�L`��C�L�ח���}Ħ�*H�{��Nl��Td��ZZ��J�1ɝXMF��=��͞>qW��J���|�v�b��4����?�m+��\�ӄ��qN���g�6pͫ�<8��d���	��p�O�J�>�7���yr����m���@�V@���괱�^?a6�"���U0��Ӿ�r8�B��o���~�:�!�HR}*ڙ����`F(��;�Mt�x ��e�E-HDc48i��f ���#�d�o���%qU�G��4��|X̜>��\��]��|ONf�_̓�(3���?5
RR�g"�gOό� )FD��X�p�V5���.��B��)��i��fL@����`����"HA� Ca!$���m�qv&ҭ,u%�;�y���H����t`�����z��GA �ms������#p�$�K�u������}Q�@;^�����
��L���b)�%y�F����כ7j6"	��3��D��>_�7����l�Hl&P�}�C8��<DS
�s,mA��?t���B1-04nR+��8m&�a�������.��yd07��7�{�~�Ƥ���1(ઃ�$�u{�\"vƶlR�+�j��[�"�T�H�l#MR�4���h??��}7xz�r�#(���J�?���I��h&�^p&�j�r-�2n���]Xs��F6םk4N�����G�k�[.��<4���z�"��@�hX�����L��@
e�b[�l6�Ā���'o9ŗtck��兰3��jY:��\^j��W������z{z��稢����N��!>��V ����݄Y4�����z�k�'R�g*S%��rw�םa3+9�͚Ϥ˫n��v���P�ރL���І6�@�Y��E^)7s�L����X��7,�<���M���<,냠�	tؒ���/�W{�R낡Q������_n���n#�3�Ac��J�#�O�Kp(��G�O.�s{3d�솺iH�w�����0x����&��4�7ݱ�Ꮿ-���R`7T%+�HD�}?3�b������g9W�kw=��]��"�v�3�@f0�0�p^�;Mw��7<=3>&��a1u�s�����e��.-e60�`��7o�Pz������y�`�i�=v��q�)����7��v���`���QU����y�t�]d��g���ѻ�rwV�!���}�'�-���lD�dƮ�\pN铭V@d��.�m0iZ+<�Hڈ�4�#]�`Њ\�{��闷��8�v�9q���(�,�������3v�ow�I��W�%@@t��K��w.r)e�v+^ߒ�#���Y�.w�e���1�������X��oK��Tgj�"��G{"p0���2)&��9�Ș�`��G�9��xW�Bk�@)�SP�<�5A8�����0�|x.���yn5��GX=����������̱_Ҋ+�ˍ��<H8!�M�G�1JC�`)�z.R��/��5���;���[�gA�mx�U>>�l�ٿ�DqW]Q�(>��F't��RUY��\_*��FF��۱��l��� �x)�;��,���%!ӟ�܂��r�$p�<�NfnJu�uC1���x�r<�c^���s��b��w@�j%%�5����B�қ�f!����̗`(E8I6I����~�3�jX���]=s��hve
��U>o�I�2��5�I�I��xqM�m���r�-����L���xBs6f���R�Os�hn@�X�Q�B����Ww���`��=,��}��|�"�S�F��b��T�K�ߺ����6�A�v�=��_�l)A�]���|
�������5p�J�~E��p�H5��(���'��o���au�~� ��}��4�֖��j������i�SG�`X5�����3����m'�V ͛�>��劺i��>�F�4�;�a�T5������ѩ��b���w��p�2j��ȝYR"W���<=���?��u�X�H�xb;y���,{��ƚ��a�c��n�n�ސj�"�c��0�����b�I�.����uUi��Ō��N#�Nx��+Wݑ��a'7�/��CŞ��i2�}���0�qa)����"�ԙ�����rn�$�_R��pڴ�Ҋug%x�uU��؟�H7s�h��G{n6�;�8��đ��x~ف0|^*�*L�d2��({4��ŁZ����q��u߯𧭺�h�N5��w�v�t��+�����Ė���7V�d�-b%>'���TV-��vY��;���7_�H�'�N����|��fG�=�9&)���.(Ih�1\�5�Fo�Q3�����ޘ��]��f�%c��D,u8~ފVe�s�ħ}p�T�8p	ֻ�,��� ?N��xo��|�c�\i�M�,��^�.�:�8wuA3O��D��֬��G@��;5�V,O!L������uE��W�),ƠS�Av�p��v��q�XeB�W��:���}������8�ȧ]̮����ה�V�~�۹XQZA�`������ڝ��F�/�D�����jB#��m�Gs�x�+r�$oQ�`�u+�88�r�N�;Q}V\$�7«��l���pQ����^��YZ\<����vJG�@l�t�h���T�Hb�f��e=�d!�M�N�6JE�[W�p@"���+�c�u��l�2V�OM��:���Օ�C�Q;�P�C�2��c2Ji�{�:ʤ���� R���f��䓕d��Ye��5]�eq����Wa�9x[�T�������Q�����/8�]}q:a]�b�候�y,|!DE����� �O�x�͑���`k(>]�����N�Snv���ʁ�.Rڽe5yMwi�2O�,VҲ�Ǌ�sn���sM���s��W��C�v�p�X���ԑ��u�a�tq�d��0�O||�͉��ل��3M��k��fJ-��*��w�cP�{VI�"d_떨��_�Wm'4��1���˔����[��]i��m�� A �x(�1t,ic;�Y���U�̳gL��m[+H�����p���{� 嬰����L��x�-�,�`�,bi@P���5�sG���z�%n�_L��tE�pHJ9?��xwTeeU�=�Tb �DZ����O�X��Ѥ��V�0NB���ZԸ\��0|�Ib���A}��a�"T{;��u�����W67��s�ҭ �"�4e\h/���h��答g�ހ�1��^��I ֫�T�?��D;�F]+=�M<�^+�c:l٢��R�)��f�䄙<�nU��\�.�C�>1�����Y�-�1QXϿ�^�ucԈ�L�/���JG��S��j�j"�&��4�?�ۋ}KN�%��RT�J��
�9h���b�R,�z��V@;�
�e�+
~=���v������CV��ў�7RR�+�,�<EU��5>0�I՝��Zq	mI���I�������V3���j�81o���ȴ��t�?�Tp����\��^�V���w���q���6s�<���ž���Ī��@U"�Z�|��_L��P.8eڲ#��t,��[Q��Ee7~ki`����Ӵ�k2�J��0v~J�}�͖����'�K/_?H��`-Y�����_g��;3S�m-ԑ��*��1𨤟���_V�$��\��� R?wa�|�%�LA��i)��d�_�Ґ">��gS�U�G�SE��IH�ozJH�˪M����'����|p.l��a��IO,��		��}E��WǙ�DX5+���n�����3�l�w[���
1V�޺AG�pՈ��3"e��nC/��]S��{&n��n2#����P1�q�y0|�c�F$��4�m|�´�R\� n�r"�+�-aS�h�d�ូ$��%�'���ǭD�&_;8FY�qv�nlE�
T��hGk��I94;�A��Y���ī8Ś�e���
ĕ�e�-�C���wX�b_��B�=���c>��g�v��LE<P(���bG�J����0/�	�6x��O�w(�9(Zz�I3�M���e�F8��~�B"�5����v�`�
�T��5��n��3�q-$��~��~�+X=�7�n�!|,s��Pqhc�N�=�(���R}���F>��������&9�]��g�����kS|_�S#����։�C�tH1�T�@/��t����OW�i�ٔ�x4�I=7O)}�޳���ٕ�����������JI��b��ww9lQ(�@"�vYH���F�D'�}ʪ��GA���'Z	և$dJ��[�=�&��}���bf�G��yf�̃>`�e��� ���l܌�L���� o��Aۺ/��i'}F��A������b.-�Aίj��D��N(nݬ�;v����;c��9\�Đ�V���6����).'��v�o��]��>0�Y  ���	���p����/�o��w�^�D����s��]H�D��x'iybX��PQj1g�ri[��a�h�;	�������3�X*�-��xX�����[��"�6�i�J)����~��f2�7]넇y�Ax�X�����孈� Y��͋#���k��o,���02~ր@5LD"^��_��\�FZôV�=������"�*.E���h�T�H�j�3(�����������B'�7��Ũ���EA��)��%���k��)0��@�)�W#����C:3��{������۞"v����{ ��-"0n� ���6�5�i�DQ��5ѡ_��5�{�"�-]
�b�'<���n�Wu]�)Jb�9����e!tai�߯���*oFWB�O�p~!���c���ŗW�HH������!�L3�T4� �}�}����Mc7�.����~�l>���(:�"��S�U�N'b�=�%$�ǋ4��ݞ@�����:P�9�w|�X⛤�v�����)>'��o�̠����{:kfX��t�\�	�7��LW�jb�5�E�Ve���Al9��q�;'j�#T�_)�u����f�Z��v�����c�'���x�L�黱��,�q�|>S��}ꝼ!
j'��2̳�/�f^�Ny��!�e�DO}�����X�����y��V X7���u4W����K����+�)YgK�C��y��O�Z0Q^��aܫJh_ba�C�l�/���y҂�P䄠*K��PV�ę�R���u�FT�pt��h��qu��Y��]_y��i����h�8)�U����&A0,���*����o�m�m'г����^q(_ ���MY/m����{Sw����م%��k3Qd��kE�J�K��������&�`G���� �!�,Mx�$f2��N�7w�,K��R8H��RY�������e�O8�o��!����e<Y�A���>Y;g�C�ie!��3,�=@{�%j��ZWV��Ȗb�<�+-�&!A�? <�0mY�}f?G�����<]�D��c�����H�[��0��n ��s��JQv����d'(y��Y����JJ�Q\&�����_�?�?q��4O���F@#�sQoe֩t�\�Y��lz�)�� ɤ5Y�R|�����s4�"�o:�Fe}c��������jI����݂ӿ��k�Ҩ��˛�֬I�p���ddn�$��Qwn�x|k�VQI��-*L�)�Ӕ��D�+j�Ǥ!�&V���>��~g�x^N|��+h�T[
Lc�{a"_4�7��t޳�.���pB8���{P�pM ���j���f��џi'm«?�����m�cw�ғI��$&����K@�r��	���|2���P�S����C�ͳ�+��K�X,�=Y��Q��������!uƖc�3�O�ݬ _\��<*p���JԨU8	b�&q��+n)O>��<�� (�&¸�u^O�� Ё�c,�m�c&41W���O�j����a��wi�'��$xVㄈ�4ƞ��庫D!LY?��U~:�＊��(ݛ^�^�=�$$@�8���t�!���6��:VM����f��-�>�.k�C��Qk�2�ʰ�x(Ad-@�NEƧ�ރ�j
ɒ	��R>��a
����.~���Fm�WT,	ŉ�zz2��T{���L�jNX�f�p�Y_#���vd�����6l��3�ޚX�Yu�?��R��hS.�2������ܓ�m�{Z�n���i�]��f�g�,�{�&+HU�{aW�%��B����09s8�_Y����Sh<]���ش��}���2��=ݮ?
C�l���A����3-�I�Ϣ�H� �����h@f�d0�Zv�ӕ&�f��gr��W�e��'9zGrm�l�����o\�xB�".!:d�$1���M�bF߫L���~Yٓ3�`�>~�G-F�iU�׿����e��H�O�i�s��^���S��k*$�<����9Z.�*ӯ�{+��$��Y���=&�T���BNO���z���$���s5d�!����+dZ
�8O��7�	%qKw�������9�9�/Ru];��8��%���K�7
�9Tq7g�%�{U��u*"V���+�`dk����,�7WlѲ�P��*O6��8^!$���-�%�M�~z�/�;�qX������{��h�5���4*�c��f,%@t�y�3�A����h0�UЉyr��R�uGy���t��\��6v�&��K$��
ۗo��^{��;"���X��֊?M/60 P���P2G�1��Kz*��d9�}����~G���1?SK��U?�^+/�� ژϿ/��h���� �q�>��sq��-���S٨D��R!�V��d XP�VY���Z7�_�ǊF�޳��p�\�O�'%$�4��pÜB�-�?��j(��dX�|��X���v�/1x��e{�{����qul(lk�&�����*��5��"z���̴�;I.���~��S��+�v>vj�S�����v(��It0�6$A�S��pc ��wA�`���Eǋ,��?"��8�\�v[�P@��|��"b _y�.F`�};��D�ʿ���L�(�ת)sچX��1����@¹�"�[�x�-E'��D����u�XN��f������ �{kF�/�,���~Nr4 Ĳ{�p�v^�����
����H��X��nOZ]��aX��o�R�s@K��~����쵝��0���x�slao=�h��}��Ý�8�=9�����3��E������F��|�mL���k�$4��K��S�������(���M�QkD'!	�o�55�㨔���o�\�.Y�`;	PO^�'�2��R�����P����ap�&���&%75��!督Tv��c��N����Ǻ�����E�,�/{(�I\܁�б�\�hf��B�� f�"0�3��}, m)���vr<Ht!��P���U���Α%US8�\�St�nv��c��&�&����O�FVHѹ"��lʐl�qlL"q�p4%���i9���=��_Ո�o�mp ����j$X6���e����Ѹ��,���O|�_�g��ez�e9ɖ���·��6��Xo���(B�b��>�ϵ�m���Ƭ�}�+�-eZ�� �G�v?aX�#��X Ϟ���r��j�d�δ"jkw�t@p��P�n�R G��M5ъ���f�`$�(Ar����"jI�RDP�3τ��]�����8@Ai_l�Ntӫ�R����v}� بu�X��IPf�!Ĭw�N�+�2��5�[(�ŭ�v��Ú��9��0��Z� �y�����-���iJ�0a�ޙD��K���iq%�wSO�Q�؅6z=�w�3K�a
�9�jE�v�Q2lvz���Ȅ��T��h�D��|0:����ۃ�����M�l��n:�)�7�����hA����US����19�V3ٲs�|�F�I���B���4׆ ���!B���ž�&��\f.Dj ���<�q�.
^��5z���
�h�FA�WEѧ=$'�ڨtF���.$���{4Z�!�ҕ�ԗ�l=k�`��WG��$�o\�$�rW&�����,�?O8��3�Ccq,^^݅��E2Af��ޞ�e���	��
��1K:��8ܻ�[$p�<�Tz�~9Y�ƫ��wX���؇�k����\e�(�������Q�%���k�;�V�h}�-�F��ǩ -}��K:���L�I�}SDlތ�̙P\�H�7T��L��W�J�kƊ2�m���^����M�al~��J�ei|���;�vD�
�(,nV�v�o�I�88%��0�Q�i�G�q�2SW��l�<\�M�;PQ	���n����8ǹC_��m�@S�UϬ�Id����ƍ+Gʝ��?z���*$x�5\i)�7#�C�pW��˛��Ecʂ�&��)���_hr��!��T3���!�H��P]��(�$Q�`�R����#�6���s�$��Nog�k�gY�W��s����$A�M��4K��>�e}/
ݼLI޼���ɞ�	C�n��#5k�A����CWɒ�le�v�j|�}�ޔ��}N�e�aԨ�j��/:E�	[c6=/�	��Db:x���͙4��Df�xn<b��.�n�xD��Mǿ���i{3����,\�Τ|Ts��{"Iy������o����Qm��{�L�}*����xI6���pZA��K��P���lAl]i����%��m�kN#WPBf��=�l����|�{.�@a��e��Af����|G'z�H���&����;D&L��|ܺf/�z]1�C�͝�2�C�V{�ۍ�ğ�}��z:kw����ц�p�\>uE��FTۘJ՗��N=W�17�����n�&H�|���^������tæ�Di��&5h:���Q9*�!E��H?f����Dd�b�Q�WHB��M�ݪ����Zxap�P��ߤ
�ݫy��V�eD� ��
d�z�ݾ|ye<e=�V����>"��If�뜶*'R3D]���Ң�Z8w���͂��tdumߣ\A$P+_�Т�ԕղ��CMp��LN�I�d�oș*�Z�$Y,��k*�(��ѱ��G�&�C�ZѺ��3#����j� !�|��zȃH����&k��<��´���l����P�����-�)J��n�
��J�^�҅T�0��p)�Xc���g�5���|����(H��k:�`]X��MVb܇b��~�4r���B__���D�����	4_�χn �r9a�M�'	��yC1��{04�JM���B�֛�Қ�� �M�� s��W3Ђ� W�(XTDc�{K��$myOwZ�~z�޴3�*��ͣ�e��*��B��GDp��>��$ME�)E���H�v�Ǵ ��WD8�L��ϳv6����A?]��!��(���|���T��?8���4g}����I�H���?�SK�H�F"Z��`-<��~/<RV��:�UT����:'̒L'��7���7�(0��߮\�k0�#�]k{���d�*�*D�K+�Y�f�$�IKߤ����N����9�L$��a�����ZC�b�۴v)	K��3�x�s�(�pR�VMO]�d{P����n�!%f���6�ա��zX�3f��������ݒmL򺏶Pj�u!t��U��Κd�m�)\:s����j�_�ۘ����uI���j\s�HP�9����,�tr!gQ��p߷�+t�����|k̡��5���rJ%�����ĮP�\�H��\��^F�`������c�U�T_S�X�L���0�;�{'f�]�[I"�%B���">9ham��k+�u�/w��!B�C�;��*%KN]������G�.1�W��`ۅQ�Oz	�����	T�*��:�M`y�w�҂<8I����0��X2������%�7�}R$������!�f �&Q��i�����/DT:� " � 2���o��Ƚ��F���ȃ������/!W���*b����=Pxխ8�!l������+�&�Ͽ�������N�e|�wI�U��ۆJ�o��� 
�1jB��/WӰ�DyH� �B_���5~^�)Ƚg쫲p���F���`�k"N��=���ϰ�!7��^�@���6S�� Ќ7��?uc�t�Iz�sQM��@L�V�B�z�Z��$fg�BV�S�/E"usWR�73�����W{�P�x�EoT)4g��s��Zn����HO�[0D�n�'+���ɗM�B4n��5}]�e ��X�l�m:��P����C(�-�����&m�V�F���w��C����,]4�n<4�/j-��݅����Z/����Uw7����\�'l��b�CvR���`�}�����>��>�p�S��٠�y�}��wnL"*��mB�
�� -�o#4��&�����Zk��|����z[�a�P���,��/��n���?�|QĔ6E�Ī^��JN��͟�5���$������0�~w���jm��j���gb'.h�~��#�����z�4$���2��5+@�U�Uň
�Hy���F�|�Dz�S8��,��<J�8�tU�Ttq��m`���H������gy��N���C�3yٖwsk��2���r�7�Q�u���M!��S��I)���9�W�mQ�H �A�ƿV&�}]�G����ߠu�S�ֺ-Pj�:� ��$זp�Vr;��'�P�%}L
�V2��}�{�W���㽖�p���P�'3�\ ��?�Ԍ����֎	�,n3|LYШ��_��34*��-W���㲙�@��7��y�r��{\�G�-q����s�wiI�=�l���5*��$z���]+N�T�]�ԡ��J҉Z�Eʊ�<�q$P��m��	;ߟ�^H<� ��ۖ|RY�./3z�	�3M۵.����}������30;��t%R*�bNt1!�=�Y�ʹ���v�di�����ߨ�|��b���ld���8�#u(3�J�c�C���WtU���-�{/���64Cx�%��r���SՄYQ�Ã2�9[ʘ5ɲ���[C���ɣ�>�#oŘ���J����"�ߕ���;�K�Zv;Ja�o��G�aaSv��(���.h�����tP�*Ӌ,���.B�B�1�j*M�{E#Ů�/À7n����a}���].Y�1�HOb���0~��5���c�c�B�<�e��F�HٌEt�~�n���\�M��7�z���0-
��,�D����c��.�;�J�� ��!��v�:x�` ս��W�j	]AުUԊ2°��[F��<�C&U~��7S]�RWg�8�B�����]�ř�Kw.}���Ɍ�q��8<��S�aP����]�Y)�P%�ȃ6����B;�?*ME�m(� nX���N ���&o�ސ�i_#@�x�Az!3�^Z
Iu���	�Ue�6^B�,B����N�A�������ʝ6����Q�#�-���lv?GM"�No�V9Zx�{4�
��s��x�����ͺ����%�@�ѣ����4m���>z�4��oI�YV���V�˿��/k���+౱[����*�b5$=�P����(doG6�h�9�Vȉ���L�Y� �� ��=V�b�{��Ip�]���U~n�F�~s��4\yE7��cdE<&Q�(��D0�ˁ!C2���M�>ۥf ��('q�`�
]��sҩ0V���,S�Af.MN�+u!�AN�~�)�T��8@벓��B#���g��5gw'��MgFr*���d�3(�b�56_BCn��Mи\��cQ�tlsi��/��_ߕ�qL�i,g.������� '�s�l*�A>UU�'�gO��@_����^�Q���1X�َ���-��#�/_aY�ץ ���p�N1�Nf�!��;f��%V��R&dW���}G�dH���b��y?�6����Ar�:q�"E�]�̓�+\�Ӯ���0>�/���1q��h?j��%�3�4�M�iwpC�MG�n¥(<��8��:tޞ�f	tZff��͹ѻU��X���n ��J��J��w�B���Ho��R+�V��e�0l 7$��мDST�a�2�N�6S�,'����l�Ǖ����F��><谑]�Q~X�����W"��@s��g�2�o�<i&*y!��6=���e�
Waȣ[���S��]Ol��E��r,���ꂎG�����4���z��㈖{+���
,�P=i��Z����W����S�e�}S�o9jb=vz�⭜�3"��.R�e���SЄh�l:}�L�Q��T�b�H��k�-姃�n`l�, JsOd�Jj��;q	�Ha����NO	��Hps��4��!Z�>�w��h�������Os��}mY^J�v�$<�ɍ{�e�(���&?H��ɱ�5#M����vN�`%kF�����̇ �g��t_C���fB��y�h�j})����WH�|�^³_����l�
����U���7�1����=�)zG��+��9����x�c{��]��:�W܄i��K�l���ζ�ęa��&����G�3��7z&�@���j������Q
N�i�Ǌ��Vj���F���Qz�}��77��{�'���ȮE͈x\�� KT���2p���DK��f4"i�w��mT�ft�	�4hp���5�~���L�ֶ�-�mqeQ��{�w�N4&����"z���BB�-).ڧ\�V{���ƪ��ҴL�Q�>x�"���o26�ȑ_W��8����#�ힲP���h������"x���<ծ�ѯ&tX�	����9��/m���,4_|�M��R���q���4 ���͒'(����qs�2�5���\n4W������U��yu,וQ
7���_��\l�Fˡ.W�����;�:���w+B����}"	w��`���ǜ� F���oP���Dù3�w;�ڽt	�P;+A;�_omw�q6:�%�:�#>M��|��<S���y_��]�4-6s��������V�p,�������-�J�}<���QZ�s�3pV�����!P a=P��Z�
T�+����a��u�Na�z��
�D��oH�$F�N�O�����c�{J���W��h�×w�W6$���N`��8���";���P?�k��_t�i8��f1��?�l���k���\�9+��� M�ݿ���Mዾb>ҍ[�F]=%�a@��R�l���'��&�(�+��T#���o��x��܆Q=�A4،b�RI���E����.����$�A)v�Z�?&_z �4�r$�Z��|��gM�$.�v���&a���=V��0�02ѹ�i���	kA:\�Nw�3C�n��a|��{$ӰŮ�h?Mm��ء��Q�ɐ�<�S=~���(hC�f���m���;4�84����9�@\��Iɟ����r�M+p8�"^	p&�R�
E] �e.�t���VF놝�6^l���]������iG,��,���F~?&G���F=�Ը�!W��B�Y2`4sz�6�QS��4 3H:_��-�W�
J��C�I�&��ߠ|i&<d��n
8|B��[l�&���4��h�VD� �����]W��5�"��,�	�^ܵI�+�Lř~4�䀭��L;�������'�c`��/��ħ�ؓ'��ߏ��kĚ���ͦ�i_�%f:�ZM�ђ�\����N?���[�2��cL�:����+�:��O��`��;���y��y����T�=vk�־/2�P5�_��8��Ds���U廎+U	2�tG�Isґ��$h�j��e�Ͽ�C(�NB��?3��{�ת�0���� `�/�z�(�R��Tj؆Jj\$�����W���i��+��<��;�f�a�m��MF&ʪvL �j/��SZ�����\b�sQ��v��,�O�q�)'
���VU&��2h�5,�KA��;�sHG}$�1�q,;j������J�=�w�\�fѡ/c8��:=^'MT��H��7wz��M1}n�su�F��dCj8�؉�F��'/q�&v�{$�l�.`
����C	&9�ʠ�F~9����ꍄ����	 �Q3篺���j{�ܥ�DN)��y5x/�����X� v�1��0y\�ݩJo���sr?�|B����gw~-Z�INV������������=-�u���;9UZu������<D���z���hD��qT*�5��������vA+v\ ��u{�奘��w�M,u	 ����[9���}ϧ�סZn;^,Y*u����Õ��ad���l��}�������nB>����"j R⿙Q�+/|�p}��`Wc�Q�Y�T�u��i:��[��w\�_;�d�)�p	����������A�,1�&�<�e�x��T�X3!T:��C�B:��|�$g��f��Ȱ�ű^�C_�C/���1�����zK�v��PsC�A2��~+/V�kg���P��E�i;כ�+(�٦�ͨ�L��6(��f�
-HDW'qbt�q\�=���KW�ݙ��<,���}g3]('�,�N����,ĳ�^L�F|���y����~���%M�A�3��(ˬ�d�̛�R�ߨ�c!�<�9�n���(�f(:�U(��-=���pRuJ���d�m 2ﻂ�.��(^���҉#�߬��Ƹ�q�B��٦H%� X��.֓�i��E�Ա�iEuSc�Cwc�A��2lZfgO�1�xO���x_�d��e�2�fx���H�V�K�Ef��`�����jʈ��8 lѰa�ȋ8[&+8���9@xd�)3��FFh@xp�s�cʇ��\���x޵53[���'�@DlRI�2�/�CGUQW�\�5�+�7�=��M�z�(�䙜,�	{~���*�T���≎3��Ǒ��(�5ת��_n�8Ý��'�yU�(���&-a�E6�W.8{%��	�A�Y۠�]c���&Dk�o�k-j�S*��JE�]!B}����Ƹ\��~%#������q���<V�����!/%a�v��U�Jf� b�X<��M����-����?Q*�p?er%�;���:(��)d����ؽ�{M� ^���e�m��P��?`c�24�7�S"��lc
�@�KӉ�ؗ �@�..�2��ر1yh�1S���P��ʗʊ��)�����F��ݞ�K�.)�J����B�f(�[|hI8�Ǩ�G����Q�ϡB�r����^��uX�iH�$��n�%-��>T%�%��t�b����Ŋ��b����g����H�2�҉@�H�mMb��|X�3.'Xb��}jY��wZ�
�«�}PdB��Jkl��@;����t��)�;�Q��Ӭ��"bJ��33akc|l�:�%w+Y��l��Y�+T��VSߣ���ߊ�d�e���j)�Q��n}�`�D5HI��ұ���j�g@��Zf+���I�
�ӟW\Ђ&F�>����
�0�U���^��1���J�"D�Խ�A/R����N�k~GH��"���p#��Wy���_X�*E% P�I^&���C���c������H��4
r�Wvm�qz1ˤ+S���l��?!�emǰ����}Q��D-|�w���T��n���UbV|��wX���~x��8o���� QZ�ߘ͚Ť&������=*���g�����	�����X+��0�a������pOxJH飅�9�t%�+~�5i#������;AO��S���Ȅ82�"�x'��~׽��Q�7g��E��B:
�>u��N�s�M9l�9P
�O��8���.Zc�@eQ[#��}���m�V���U�U!�	��"N�r��Λ�ԩ.�2T}�;�Ƽ����) ���1"n�-�˶jߠ�
�G|��xZJ�rt���ط�M�$۩�EG�'�)�ZK0Z�� +�$v5�����-Zbo~$FGE(5�_0��b{����w�Ǔa�8���g�����ad�u=b?��;
$Xg���ğ��ޮ�l���-�1�W��ER[[�)��|�d�������M8��W�ҡixW�?��ۨm��I�me$Ds���pa�m �z8?^��}����N�?��Xه�)7���1�_�'	�'�	(c��}I!G@W-�B[�/�V��V���L��� R�&��)i��-%D��WjFX
d�	,6�P���M��bt�y]t�#�X��!�nž#>7s*����ͳ.j�"F�m�~l`7�Z��p?%�֪Z�DEМ��"<���i�AL�Y�l��x�zS��1L37�D �\�9�#���M6E�H���Vxe?�
 �|�u�	��mغ@��@	!��t�C��X�Z!���J��L.S���Z��b�ƤZ9���*�
z<^�������;1A�ͽ1�Pp��/|?l���e*�H�o�D�����v�&͔��Es���}�!�������)�J�}f�O�Ӿlf �5fJ}��ml�K�e]Yӷ8��Bz�U$#܂�6%���?Nie_������/�����%��q$pG��pgȝ��7�n���!͉w���eeM���"��|�x����k�} _��^�7ܕ�!���zB?W@�6�?=�Չ�\�9�U���2�����f7ma���b=�%�������/+D��T���D�)oP8z�c�LlE�����v�G	*B���+/��8���
#g,YG����9Z����}Г�	
.���?W�r6Ц8b"o�w���+!�ՅM���wc�N�p��x�1V�f�nrM��b̬��A���G�h���J�G;3�E@^�s��E�˂:8�4���������g���)V8�{Fg=UV)\��~����@R�c�i	����BxN(�4�;'�9���t}�
B��,�K���P�(��uj,��m�2y�����}u�[\����4�F�]�p����v��_d�3Eo!͓�s���]��&�u���K>L��n���	S,�����d�V��i�Kn�?��1S�S����6avFṢ|c�δJ7���`C��h�ű௕)�GJ��W��N�:z?Vb���U�� �W�M�F����wB��5�hF���g���s���8{��`֚����#��	r�utWķ鍄K^�$F����Z-�lz=Go2��Z[��S�%�Q�y��v���x}aRN_u�)G�~�fJ����#qAZ��J��hQ���m�����6R(�\���9��ً��H�J���w��:O��o��dƵ�]f`N�H7����\W���+��Tj� ��Ҳ��͕��<������k6e�zP��K=�=
��n�!���`�G7�?i`<~g�|�:38������"c�[M���ك�� = ����_v&>Og�@�C�l6R�YY#����^�ʹwM�hq�4�$�e;�Yv^
��fOëo�9~�u�����ñ�.o~!3��W�|��j`��x� ?�z���c��˦��Y�;�����o̽`9i�M36e�
M��:Ez�Z��X̞��l���j�� ��iR ���3����'~����Ҭ��F�*9+�~1��Z���_���䳴��M�1�F��JW͟��TZŝ�0QG����d�]����Y��Ob����܏%:j�^E�dc):�R�錸>\�Ѵ$h�@�[Y&=�4x#,�,w)L5;���`��E�;Nbi0M9L�<�1���xm��������r��J��-�U�E8�i��!k�<�n0�6�g܊�B�Zlۢ˼?".�!]��<k��˗x혳b����A.�.�z/��� ����&ah����?��yZ�WZ�I#VN)���v�,������]�B�׼5��$	�ͷ`]�{G��J�1��^���Q+U�R���2x<�Ę|E�N�ݴ���Ww��ft߼D`�SH@+v�A��{N*�!gr���5t�?"j�>�ok�[P���K�I���Ӎ0
��>x���adM�^�U�'N��獩��HN0�>�W���m.��cx5�09'��R!�)4�����ɧ�co� ���}D�0���]>9��[��C�46&d���V�Cm�߼Y
6ݟ�2��~-�zI�BhSq�4s�P���+v���r=1����Ĭk�]��մ���'� �,��^�|}�T���M>��0�ʀ�gxVMQ؜�\����	d�o�~���(���'m�^$��*�����+�D넪� x��F��{:��c��>��	�ٵt��U�d�8�|Pk@��������`����Ί�]�hC��X�o_��Z�V_t��C�ݗ�pT����a�c0�F{D��hPLw�,�d���K���u#ù�p�Eۿ�B�8�����^��-<�"������:���h������Ş�q ���v-OKu0p0nľ.��"
A����-�M@�Q-�$�Z<�m(y"> ��5�k�2�ܣ.-�D��6�_�cR�~�ڱ�MY�sK��G#>��=J�L��'Ks)��_%�Z=$�l�0�\4��|_=^ˋ��ڒF/~�[Տ0
�P�N��tf~b�����!_��F�C��Z��|sRL�:�*i���#��gg��!=�Q�S��R�zU�*��H�]% =ݷ;(CԌc��B��X�f�O�'�4{7+8j�b�Xh���<3�&�3".�� i��UoW��56R��_�\�7ϪJ� ��1=��|�]�G�ֹ�K���a>����'�G<o���h�Zi��eƀ�L��h�mSY�]{��.�5�?��[ک�����Mx<� ��O��xp���4U�z2Bm��4"F���A�R�`bQ���8�Ze��X���f�Iu��/r��.L���@�j��(zkX��1�O�]���!�e�?�>q[c�ѧ?� �9W�tL�3�Ĳۀs3�	P �G���Y������%�7���1�	�m��A�cy����'n��Q����4�ǂ��� 	�R���%�������b��SC~���-+��?|U&�0P� MꟋ��}׶�س�!�����`�-w?�a�����.¥"�(3ϦtG1�h��{`��A3�Bǂ��H$�mD�P)<XM�R�ZN�{��.�Rp1�~�R>�|�
�9b|Q��cͨ#��a�ԇ5��Zu�Ha�p���(n"v؟Y.>3��;H���_���-���9�y���/�*���ڗ�}��^?�Ҿ�U�Qᅊf��?�vd��8/P�"�ܵo�*ND��v�����BA����.�g;`��89��|@��	�MKYi+��B
�Fz�w�J�II܍U�	G���t�������
��V���r�\Tj�b���n8I��m����ޤk#a[cs?θ�}֍9V:O����f�B�����h��Zj~�^oB��/�@JL��O:�O��P��~��B`�g���f�5~��1	�������=�B��
~��u����.7���e;�D%�,���F��a��0^w9�d1�`�����Ï�ԨW�<n����#
�Ù��[i���,�R2ь4��T����9�� Ƒ;	����E-��F��R.m��Y5�\�jÈ�T�Qdh?Y�	G�r��9�Q �D�=G2�d8?�K��+lyoE�~W��!^W�jb�⾡E�6T��i�Ҩ��JP��4�ܔ�i� 	��؃s$LE��"��DaI��A�����S���`3+�{:���Z5O��#*�H�Ll�n��݁��fPi��W��k�����U\&��|F�RN��DB�2Zf�:�<S�5m,�Am�hh
 �^Nd���x�.㋘ֳ;ӏ�C�"}�бo�C��d=�Pb�ٮ� ��qvd���G�Q��*j���c~)E���
T���6���j���#P�w��[�?)���>\���@J��p�}��t$?ͤ��-���R�,��l̿���Q��g}��\��A�ď�����F�㨑���C�����oL�H��˷�\�bU#�/���F���9�/A�?�8�;?�j��={{P��:p/a���R۰�`���� id�������U�I��{$a���Y�E��~�p ��T��u0��߫��w����V]x�v��Q�5kc��9�L֢���γA��S���<{\U����,1u0��Ks���bi���Mt�`1��
Y��p
�����C�Z�y��O�'H��Nl��./(��nҗ��Zp�����
���t��p�+a���9H`4���Сg�ߓ;��r�mcGP䣪I���
� �P�a;�;�]z��l�SQ�t��x*�~�����A_Ϛ`�H�{AR��t&g�#��h��2<9ق'U��I`�
%D&G��4{2��M�X��T�8F���;Ȟ*^�bY�7/� �8Y�~�EC��W�:�ɠk�q���I^���S��n\A&����VPzl�X��Vم�&2v�;�֘�[���{Ջ���o��x��|߸��V�I�kl�}�|6�̲���'Y����QB�j~Cm&ޖ��2�e��nZ"<f�,t�8����j5I�����u�� ]����� +�u<D	��n<<n��#c�N+�������V#!������T{��ᾞ���P�:�D�z�n(hr>C"R·(��Gl�v2���ޭ1���ύ�Ǆ���q�ə2���8A�s�5%oZ0/v���Ί�#WO8>&$�!̡2���il�bϭ��VQ�=��&t&﹟6˼�>a��s��p}����S.�R2�"A��}P^� ������l9H�n��j�!����݉�[� ���@��@ ����n)A%�p��	ዹF������.\`�H&@#N�`9�P�灋�$Ó�ԓ�ڒ�ά�W��J�����öp<���4{��t9��r��y��tB�M⎎�[By׵�������Ť�D��sܪ�<1�_b��A"���gmG��{�$��8�R�g��HRb��Q_+��dQ���;w8<�^e"!)�ǵ.�^%�Hn��pT�'*�%|�W�tQ��6�1]�pD���2�W�䡢6+뇸ERV��t�Ȕ���R�/�6f�jB�Gu��I,���7��P>�s!:&25�@��P�O�9���4�h����� �j�v�^Fٗ<R}�wH+�<��K1`������~K�݈��c�W	d��� ��	Y��u����1��R�����rN^��)\���Dm�Y��ά��n,0r�C��j�'I�[��%����3���ܣU.'�if�G��k>�eU��@��O@����0Y�j�`$&�_�^�|��j�m#\k�(���Th契��d��l�è��g�p� �""V|����Ϙۺ,��49��{����_��Q/��5��9=1Pղ-�(�l,Յ��d'wx��2�Ί���r�ޠx�X��eGbz"��%Ui����O���l�7��HƔz��k�:�
��Ts�G1�Xix|0�#�IX�9B���hv�<vPK�5�a���Sfҿ �vZn�*�x�yws��.�X�,_�U6Yq�!>���Fճ���A`rZ���n��&gH��(j_Q���H2��άV��1	���ָ:��a9!'Q'_g'E~�z%������
���{eM�2b���O����T�g{i�U���mԴ4��G�#G���A����L�Go�]�.Je���#�9�1���c^�h��l����}� ��j���FB��7fo�鷒��O^=�c,
[Р�ӨA�@ۺF��Ô.�ӿ	|��D�w�H��vq���2��#�x��?�X*��F .�(�8P ��(�8�<�t�$�E���h�U�4�J<̰G
��f��ͼa�$W옵�ϓ��Y�jǣ��;a�t��Ζ�C87��� �� ��4���%\7�g[��k��Ǒ m	�����tl�٢N�5(�߼9m|���{��˯)�<;����dSG�ڂ�N9�� 8�~=&	���j��6_����<����]:8�N����_�yt��p�S����y�KhѾ� �\�N]^�6�#Ӿ\ӛ��G{I�
���L��zώ׃e@	�L���2�S�x^�FÅQ�.O����ټ�{{�%���ܹ���m"¬��R�UT�h��/�ӊ�����eCd�6�;v�����U�~~fy�8Q��w��x ���ҥ�ɍ5�Fz���ȅ@)��x��y1��љ�to��w�p7)����wj��3��6����/yv�A���'���?Ba0b:R��JJ����P���GܘҎr�g`|�;�S[�_\H�_#�1d'^���DE�A��$@D�d�܃!&bj�j{���v�Lut�t���1�*]ћ���ת�݂�R҆69��U��&���,�����--�=U�W�Iq�� 4g"�UW8��祠�<A�9��3W�ޜk�>��-�΢��K����ٗXؙ&j�t���'�U֬�5���Ji��hD*�vM@�z�J�;���6 ��*nl	t�uC�W� �9Xg[�.�.�G9�~ǈpԧ�0�}���US$�BUA ��Bm�8�@���3���
�����venUs�
b�8 ��+r]�A�JtrH�	�Ƚ��c;b���S~��_:�j��Nܪ�M����Kg[�E�?�{֍��l(93��h�(��=�� ����2H�2�3W1��ɻlF]`�r���K=�1m~�W|���0[,ԇ�AA����$J�A/�	�����퓠��7c�}\����p�5l������ADִE�E�#_f�7H��if_�Dm[���>Hs���i��x�6_`�fJ�����G��M@�^�	��R9�o�/�B�~Т��z�����
J������!��P*+�d��)��\nqa���q��v�^�}d���'@	�3�y�?~���YvޒUIy���_t�[Y�څ=Bӫ3hU��5^����	���ɑ��,��[���J�LNv��&���W�ϨB��C���G�N�`@s3�Y�@s%�z˲!�s.-��n��7ʹzɚ����v�a�Ҷ�Ŷ=���+4�)5�"���ۧ��S��r�n�qdj��l��z��<0�b(p��M�#j��`�`�;v�Ǣ����4ĭ#�ډ3T�y:��s���ky2G���� e�V.�
^{IF�@]��n�ՙ���g������][V��=td�9\J.Z}ċ<x��G�������G�Lf�p�y�|�|~�ҘI����>$9:��!l!�� �`�>bL��x-H-;�q�zP�66��u���~��-���� �{z9�rXCo�#�2*]���?���|N��9�L56��/T5������d�~�L����Wuņ�
�a1�U�]0~+��S��L�R�9#jD��MBqT�� |�\V���[�3$�0S�I����=��µ��97>aԬ�q�+d���qѬ��,��?pk���t��; -�"Hݻ��f^|�,ו�E�fO��Sᢍ�m��a�Nu�4���iV�1,�7N>�����1| m�|�6M��f�j6��.����+�v檶���P�FA��u����B��B��2Dť�.�˥��Bh�㱩���I*t��Ti����́�`�*�f���0�T$�M�IL��j����ۇ B��~&=S���B�\6����! ض�q��D�6tr�À���L����u�Ҹ(���h��0&|)�g�7fsÈ�%�j�^��z��ڍ�#  ?��2V@�����M�|QU�y�f���	a�5�\L`ޣW4��ϓ�������� ��o�|���� ��I`e���SZ��w�!�u�� 4*]�;��s��К:E1�V ���,lq�c�c��/�dRC��_��̍)1��É�?�	R���*FF��������l�N�T��SV:���jݷ)CK�Iv����WWc}-SQE�c�z���jO�ߎ�Q��d`x�I&R�4o�,����z���
�Dzb �|Yl2N��Ju��\WUҨÂ�l�eH�R=�>�DwHĆ�*M߻��.���WE�JrJ3��J�HS�������༜J��j�i8�x�P,>�����.�kڒ�fY���0�f-���u�Mjm�%t6p��4��{}�t'���'�v�v������U�1�Ny��_� �"�8�G�'LⱮ����N��D��bxМ?RIf��"�YY���
�o�U}���a�@�Ob�;@j}��SAJ�*�,M/�N�X'�<�
ݦ��U�GB��:��vl�[�*��j��a����X�"G���J��L-I���j���m�+��wY+�=���
E˂Mͱɽ[gNW��ַ[���:.N�ȷ�o���X` I��	>@���g���;n�!.�M� �𥇝X]
r�+3�^M���7�\����Vp'{i���,A'&k��Td���=B(��$��U�ǹ���-K�W�H��ᕡ�a+�	�0w5���Wv�{bxN�T2�=�f�����8���U��BT2]��0�uίE&���N=�s��,�ُSv��	���,�*�ǖ�%�Dx3a�����'��*ힸ/���3^r���f�4�k-�{����1�ee�%�ݔ�&.��b��D�#�&߾+��@��58���r6łt�Rܥ������2��RY�g7�tS��fW�Q��\+w|K�y�i�F��>85�h��ךZoҟ!p`��+8��ɗ�u���,FϷ�P�H��9���^ByJ�e+#����]��6q��6c3h@6����0�}����(<ɭJ&0��᱈�Z�\���o]��\+(�j�!�O�aV������W: YSN_)�oL��lp�}�������� ̮Q��B�ˉ3�i�K!"wo�]�	�tm�+����	X.j'ㅵ�rS褴�)�d�{x�CR=�om��/�p�:#���pC8h�Ԯ�K��p����ݱ��da�0�ے��{�����)��7�X�Dɍ��:Vu,����:����J�H��ur��Q	����D8$�	����1rH8H�#�f�y���}1�ָ2����kp"?��)Egdx����u�Bޙf��*��I_����k�n�P�v�"�;�~��yX��))��b�g�ݡ�./�d鈰��k���4�(ռ)a
#�zf�kj�oږ^���(x�����S�����љw[�m9278 6�!GhSY�wUK��e�X�wS6ꑛ�x�yVi���ݕf��<s�@�&�&�p:������xE"��b���S��5J$@3,
�a��s��.m�����~��-1t��(?H�����e�r5@���V���!L6�^ř�Al�m�Bf�#X����6�������=F.CF�4kw2���r��Ĕ����^��M��-ѵ��s���O0�(i�����@@�*Jh/�y��2s�y��uUu���3��K~��R��%64P��oJYv�21�w-�f-ڱn���@M���]��T�0ʉ��vW��� *| �଩|��/pjoR"i7���P���S��Q�R>c�I�SU����z��q" �J��4��g�R+���,Ǖ "*��c�����1�3�]�c��W���R�Ƽ��Pe�p�^����K
����p���IW��)�G���7@�WI�T���M*��]�2��K�µ�'����p�
���!p�;Xa����i�T:�)�+�	�`��*]��syze�X'1�*wJ��K�����������BLoc��?��E��mP\����%�}���&"Tޤ��^�q�gϨ9���޼���@��_L��a�x�u�X��χ�� :T�'ȩr��"�������������O�n���aC��tO��j�  �t
u��ڝ�\>~�.�&e��#� �"\G����A��vY�5� �?��O���p�?�C��t��x��o5XM�c�r4�Y7��e�^�9s�%t�c/�6�\��)`��b�Ʒ��uT@��F1;��%[�w����=�¿E�4��o�j�$�����	��{��Y6��5_����l<��O�؞�4�H0o� '_��ܺ3� q�7;��{e��"�x�>�#��~��w�̸҅���]p��
9q�Ϛ;?�g6���H�y��i� ���{�qC����������T��?�"�el��(M�&�u��[ѫ>ɸ�8�f�����P�$��B���d�Pl�"�>��Jk;	�]�;fu����j&�Dr�׻��i��D	N�JѺ�[�z+�<�ـ��m7W�k.!�&�v�i(�Έ���7�{9��[����ª�SE#Z�N�#�lvҝÕ��3�t�����rc�,�����2��O9�@p�~����Ŧ���3aA�%�#�>��58a���7s�'�W9��`8������R���E�:?�d���?Q��M�f�����tH����K�.i�la��Ʀ��͜�hų���f��_�,Qu낣���p��*���1�N���N$���T��&#%B'�\\g�����>ŧRF�8i K�-����+��@��=�d.��3W��(G�Y&�6�"Tz����c���$3�� G:�ۻ�������1�i����1��*�#�?��s��HF��3Mr�{s+�1�'^&d�.	��)�)�Zp=�2��?������ʵd���^���L�R�9�8��+��������T�_�m���4s��{��Q>�I^�F�q�9���N���[��;��U̽�oX���W����:�b�=�ك�@�
����b�엨O�����;:��2i��awo{������� �u������RԮ\��.��Y v}�iRPܼ�`b���B���,�u�]+�t�-b�Ԯ�G�e�hr5���O>�n��Ђơ�y%B���բII�V�Pz���u����� �|~����Vf_[��\D��_¤ R֫�M���\�u]L��]Ɇ�K��x�f4��e}��#���~Eo��u+;I�UX�F���T �y���tا4���6���p磖��Y�Db?�tw�i�Qc��"ڒ\Jd��@�N���.53Ԛ@
'��}�XRx獤������GӠ�oe1��O_��n����~�O�z["�F��D%��m�AF�2 (�3����ev�"�jG'utt*�����s����l��~��O�v�T{������e#
4���eM�_&���W+�Nu���]T��t��b8>�`0i�ͧ]��[���8�Y�f.��K���N�Xԓ��!�jr��k	�}ܥc��^�u�h�b�#Y���H`���F�Hq�H��%��z#�CT-Ӧ��(�B�)�Y)p���]�# *9�Ժ�2�A�M�g�B�c�<T���$?���,�fee� pf��D_�(p6u�;�k%�9�&=q�>����+ǏW�B� ��%��{|�K�
�������\.�J��&�Ԉ?n5SJK��{���l�mcr*��]#�~�3;ڕ���O{�m�`6?bP���Z^B��g��>��.����=��W|G)4h�@=3r֪��k��˲<��j��k$�.��~25�7~���:�瀬�N�΢�	��H%x�Ǩ����N��\��
sq�z7z/�e�#b�Z�P^}�w~ѭ�7"�sp�X���5�L����ѣ�˴%��#��t	O��}n(�|mZ�ɇ�����a��7uX�^����/p��9�a�T=5S�Ж��όg)�(�k۷c�Vc,�1��7��?�<�ANlNy�a�����W�n8�5����$�$�]n&���ihp�U�0۔�^Ã�B:�8nH�?6z;�� �2v��B�/�j0&@�2�d�V&�}J��T��]�l\v�1 �#�O%xs?�ʧꎳ�o~$.'��c/3�TQ=��ˈ9Fq�ld(c͘�!Ds]]�d].rI����d�dR��O�cv^�Q����q<郵ځ���Q�4]�L)ƨ-�~=��Ca�Ы^�s��׸.�;q$�@��%���k��b�H�8���fܡڅb� ����ioO�� �Zt�k憑M۾�.owL+#��7�Jɉ�,=�M�����2����-�>��j�D�P/}
����P�/���H�T�G��3{R#�L�%�l6i�"ʄ�k<'����B���WuD��U�`�&�"#�c(�Wk^�]4��_�]�X�:�Δĝ��`I!�bk�/ԣk����sQ-ؙ$B��K��ߍ.A\!v�ί(��"�ss ���g�I��btTT���ST�p��)a�詰Z�X��l�yU5�<��TW��h��#M�XT�˓�,������S�<5b҅��P����T��T��x�I<>82��*���
e�i޺�	Pn>fF+K��f�D�+�rmui���2$!�y��O���.�ta��oU,�m(���d��3��G�C��GR�0�����Q��F	�`y~]�Teߞ ���{ �Ո�nL!F���:Kgt�^�6�e�.���GEw-nr��/��H�P�^� ��������o��ɤ���Ӂ4������}rP��d�ÑѺ~�������^�����Od#R��N<TC�feu&��VYpe�T���@���.��*�ې\�N�Iʅ��fs��t���k�-�y���k�	A�^?m��D;c���]���&�����%xں�L;�'q����c�Z���� �<Ns�]�c\��Ћ+�B�E�ǩX�g_��QG;8��w!e{R�y
�*B���i/�pR����C�|e4�Э�� `�TS�G���I�t"+�z�b�m@�����4�Y�JrV 2i�z�Z��uV�W
x�?���o�Zn{ڥ��^�u
X,5T�?��JGӸ�;x����8�{����9�V�z>`�ȩdjq�ĳN,���V�P�H��Z��[��@�p 8Z���rxn>���-�ȼ����vZvq'��Fq��gh�8��<)3t�f�ٛ)��Le��A�ǢHF 1m'������/���ng��������PWh$<)�@b`��9��'��Hؓ���a`�
w�^ b(�	�,{�a�Mp�"iZl���뿚�|��V�х���9G{<A9M��ka%��*���^�.�3��k�sx6�g����]����+����6P�T�Fa�k��Z�A�dd���Kq�.���>�,��G�h�G���w4B�Q��YWh����^���e'�OA�0<:5�����v����?�My��|'�M-/������+ntv���&W�[Xn�E17~v*��䨊 ą�NŨP �g3�B�&ڶ�R��{�ސmO�5têo�E �5����� ��U&���PE��|J
�J
�{�+�����}��D3��aX?�y�M@����4ecdb��ʙ����8��,laà^�H��{��@�/��|��B�)����R�V#}7�ͬc(�{8���_��uH)�����F0~#�j2'H���#)�pK	�W�	�J:R\//QQ����p���(�E������H�� �&xSR�=y������|
���S�'h���ÙO��96Ճ:m9�W��-y.+o�6��l�8���6��ʇ��\�GQPa�@�I�(�+�<ljF���	WӞ
E|�[�܍��2�ŶC�:Sun�!��eғ5Z�jn<x�t�r��s`�~n��R_۝+���}P S���7<�&#ѷ�<�a���R����R�����=�7{K2ȿ-��X��*m��ux��K�]D�|4K3��N#�i��
J�s�W1`�h���OM	�t/�lN+�׽��U��Rj�#�k�g(}�g&�f���W�ڇ�u�-��!	Ac:ƓQ��>5("��G�� ��c,%k�\�@3nDS���ç�\��al']2U�dS��[�s>.���ȧ@��������^W�3	���}9��ph�Us�j���Z$�_�Վ���-؞V@���V�
�P�=�]I� �%)����eA��<&밳̀��Aw�Y��S"*��E*�d�.x�YZ
A۞��B{��i֯�C_��=��-;��'���j,�w^�v��<2�ao��Z/{����'+42�OS�[cu'�3��;_��ev$9`����S|���e����9w��0d��1�ӡ�Qߖ�5:�(�½0��1�ㆋ�;�~5&ʼO}~9obyJy��3 
��H!�����2��K\��B�}�G]��A����e]!T����d8&h�σi�b�ys�n�ʏ��7DYiNΜa���|�f�7�#���_�(Wv_/�}�4���&�?V�7�4����,�󔧙����Q��J�o�y"��A���-�tT���h�ڏY�'R�8��%m�	`Kh������FU'x����- Ը��Zd�M�~/;R�Hv��e$6b���F�t�a������Q|���f]m���XU8�c�-�C+�O/�YNo��!)�-�모(������N�$ �Lm�sKo�#�/7(C�UJ�T{7�&��
X�'���gAu��2:�o�X��ǿ�V���c]dLP�,�j�Q>T,U�_�v2�oj� �y[a�A����~I �Z4�t��D�5�p� ߜ!����CŮ�IT��w��xJ������<�0�H�')i#�
k�v6$$6��bt3T;t�x}wr[�}����m;aDc�	a�ɍ���6��(o��Z�]_�텂��c�c������_�*��f�``<�R�e�� �aƹI��D�G����Pa���<=�����чީrs�B�x9�A�9�A��p��P�~�A�_Â��m�OW?����r@B�;��e`�8���}>�6?�34�ݗ+##_�:@/`�N ;-[��Aǃ�t�pḓf��5W�wab�|E�CsV@�3�%�3��횒���D�Z&�y\=��$7���^�ʂHJ���0��5�2���C�e$]�E9��=���w�=M��`��%�ӱy.V�7d�4P��6�����K�+�ee]q�'��(���wg�E�{��-)����hR��u���~ۈ��0O<�|U�t��KZi���KBqgf�����t�l�޻x���V���~�#�0��܉�n�:^��7 ����]�'�8�����0��W�U�9n7b=����7<��� �)+��ǴHF�F1#=�ߵ̵�1f�/F�kD�x92�f�ΐ|>�K�����1�/�������dJ�v�F�e6�`����N����:[h �����ל��	2׃A����B�Z�)��֑��Ba��ėW�c�����k�2'���6�EAzv��-��Ѩ{���&E��ů]�HD�tގ�*�Y^���Ɗ�yp�/ �;�ؚ0�9H� �[_}�
�J�`����R<
UAM�6�K$�*����b�["h��gz�{^�q��2rnfpX�֫��=K�(���I��}�G{�v��N�n��� fF���]��pk��j�����.�3��M�;u*�峻��C����D��B�|��ֹ�o�@�m~�8���V؄E/���j��� g�����}n'��·��p
���?X�Ԧ%�b_X�KK����ٍb��JO��T�vԁQx`�𐏠�i�{�o�<�C^������Q&�#��栘����]�;��h�His]x�=jݙ��RJW��W{�5<�J�.�xӎ�����;R�ߘ��-�9������g{���2�����S�'�������.�Q�Q:d�A�Χ)%�y,�� Yî^�ы���V���o'����ċE��_�"-�SL�W#��]���R4��R��� ¾�|��m����r胕�����?����Y~��\�H��qH�D���[���J\~�T�����NMW��0���
��^�%B��*�F�ݣ��%�:��l�I�XԓA��7C�Xt��*��щ4�-%Ӭ�;6}v�d��WF=<R�}o�����5`��a�R���A_���� ���rUbI���8pz�o���
�ִ�:T�9g�E<g�m��*f���E�J~i�^���j�o���:{�?ޞ~hU]O<'d+���*�چ:���[g�ܶ�빂��;F�?
�,�����ʑ�؉sE�{���q��a�j'F<Q����,J���_a�3��Zx�KC���K?]Q�V}��È�΂x�����"��U��{�*�,6����e�ːI#S��D������cL��P ���P��l0)>Afp�G���^%*t��fg�E2ce�!���)8`/Cz���5L�d��ʢ������Q2�i'Ք"+0_����-����{Z]����⫺��&�g���!�SȈ�@�[t�@���-i��B+W�竤�Ҭu���{.n�2��+y�6�h�W�䝼xl ϲ���4��8�P�4���}��!���dk�W��ZJ�7qm��60z�H;�o����Aq/���Q��ik�_�?��I}��I�?^|��$VHP�3�����Ǒ���	�p��x�4m�eْ�uW A�r͚�n3�\E�,8��S�c�������p$Y
{P:mf"�+d�3y��N��0�I£�0E]�?�S���z|g�>T(�h�n�_���$E��
lm��vq3��^�R=.qؚ�q�d7�|��|�36��'�*���i����-)��>I�������^�/[�I�:@bSnaQ%��(|�Kв&S(0g� L8>� ���L����L5��+����{}(�$gE1�}���)�L!�۹��
��2i#�#Y�?���Ȃ������y7��'�;�������F}H��bB�$�@ԥ#�� ՞���ٺ�gp4�$D0C�nHƶhjw�4������:����ݝ�8�F]2��6cr��J3X_�9cF��"�����TG����-��Hi]�&�;�D��v-l�Fٗ�L}�֋?�HV�lH�+j|۩LZ��U�%�aT_0����t~�:-}�����>�bwiO7*�:��-��1Wg.��r���ގ�~S<T��J�M��I��5p�,w������r�����Zpd��Ȃd�6���s'ѕ2���۟��?�F��^%5��_'ϒ��2�hh	e+��2~1�X��W*��@N�1���L�@Z,Lt�q
ZU��8��+���-���*v���	
��a��+䂝_�`��[�P�Q�J���t�k{E���3��@C�r ���}	r�l��HJ��Ԇـ��4����BF�c�}��e��q"�f�)�����W�5�>B���,[)�g�����;�Ӿ����e����FzŖ�V���xD*�U����`3�';�a�� �R��~⾵k�f�ӭ�C��|qh���2�%]����Q̣^�%�M���� �w�.Z�v]Y��GwC���e�����Fy�i�����GS�w2�뺺�吣y���<��&|�V�Д0�jE�BF���
�ɓ���%�����ޏ�nܥ͆8�ħ�E.�O�*�'��Z�{T�p#�.:�GWu���C���"噇w=dA�kw��ɸ��-=�U�����՜'�(\%ꯒ&R��ڱ��֖r_ћc&�gk�����*���j��o1�bc�a�fkL�4)��ٗ��Gk"���E���g�o�]5����0`]�p[����c�  ���L�C9��2`�;�>,��%e#��f�R0s�(��-�t��]��aB�3qVͫ�����Ō��a5F����e��1^k�m�z{6�?o�dN���$�>�/�8�KЃ)2Z���C_kR�ݡ^zi��F� ��� _[�o*��K�g��v��Q"�-P/'�C�)ؚmΧV���5=(!��SW� ��ѳa�8N_.��o�$bTdR>4�����PJ�ox������;��B�^˞��B���`-E`V�|+����Kג��8C3����Z�)���p9U�x�핬��8�H�Yu�fD����n�ԚXN��2}�p��X���-����c2$SeX������\����T:hug�2�ǶW��7��X��z��^T@'�iX9HP���@�_�%I�x�ޕOg��WJr���v��^�/��\�oz��0�K�¦�����D����|X|Bs|%Jɤ�<8ˑ����9����� �G<��F�ߞbR:�%r��SA�E�s�L K�����0�s���x|Iq��sL��dF��+�������L��mu�HN�^k��&�%�	~Y��Ӵ�Hx�zi.�"!��h9�f��" mL�ںz͹�ځ���$J��������ij�J�Q'Vlz�k6�~���ӱ�w-B��q���A�b����Rř�T�Ɣv�&6��G��#����w3~n�����9r�L�Q ���BGrw�=���#$ ���O�\�tؒ����=���ʣ^ 1�@�\�1	�D���mJ�p�4e�ն- �c��f~Pcf��^dBz��wJ��K�mV�w��ȗ�jE��>0�ȝ�y�90q�SZ�a�F��y�L'�s4�B~�0�F�����D��_O�9���;0� U�6��vVc���a��t;-Y�{���^���GFd���w�v�rh�'������-���D;�>��r;5"�9Y�5j�R5G�]X����+N�����6�,n�ޝ�ކ����1v̬��C.`I�B
o�N�ѕ�jRTeI�gK'cm��q�Sb"���"�Ӭ|��26��x�&��)R3��N<f�[��'�� b8�L�.b\�k�n�c�e�a��/�;���m�d�R�/|Y�u�%�'k��.G!�~@����9jM��-;�$��\s��boM��*��^,5�$j%S��ǹBf���Heױ������~��5P�f��SV�d7 mu���Gm̜��*(����3��7	���@@B��`���;\k&Brz����-�E�?�P6(V�CE�ٖ����h?��9ʩkᆪ8k`^�!�X�6�p���aÉ����pHBu'�ԵO��:	$pW�9nlWcp�(����Q��Ͷc��c���G}Tb��-i�EN����
�?�Qu7;�o�+�����K���BgZ�|�x]ahoצs��B9�=�B@������Ktpq��/��/�~ {���b�/0�a������)��W�2��}]V9�S�S�S������ɪxq���U]Ԕ���G{&P�8h{�����'Z���ߣ��*/V��;*���ݧ&�T��싿r���N�>�����t&qb�f9�W��EԤU��̅Z���ԯ,MAְK��<M.���ɳ�&�Q��"�+����#����b�J�2wb����,�GOt,8}��J"�鸶��}!�H��j.Y�_f��E�ʬ��R�7�C�-����z=����l{�����幜[4��
k��^A�72Q`��;S47��X��+���g� �}�{�ĵfMYYվ`��u�(.�u���
Evw�8��7���j�wCOӡ$���im�"���j)3�>P��vh���|��0�8�tN����H �Bmx��2'��������-9.�^��g�,�"ܔ񓱴��Jc���r�ҶT�0C]n�w�S��#��V�[%Bg齧P�K�C�]£Kw��Q'Ո�K�����!��򯜒���H�f$EKG䎠N�'�猋��=�5���%���3����"����/|�� ,�����1oxa-r��ff:T���_Ki���!�{h�|6�+$mw�c���+�ma�Ա)V��U	�Q^EM*�{2*���Fr�2�3c.}��O�!Y��5���Qu���-p%��bp�->�z�y��E�"<)�]'�΄)�S��ռf��铢H$���u��	�W��\`�J���	������k*_�Ŕ�8�1S���>P���?�IM��0J�$��!�����r��\��8�a���e@N���K�Y+��)�|��dutz��7���"UMTM�x\����`[�Mp57K!Az�j�)��nWn�<���G�9S��j�_�
y���*�P)�(ޢ�J���qqQ	�/Ė4�8K?��7�'Q��>o����bD��);>���^�6�+�-��ݫ��ٖ5ˎۨ�3���3 �Q��Ux����a�Y�����*E����״ؗ(H����ŗ�=����Um/����Y���Al�N�&���]���$�?Wl��0�j�3[����K��}�@KJ2��O&Ϛ���P�����vBW%]Hĸi��@��d�s+��[�Ո��w���f�?BQ���Ӊ7��,��1�!��r�k���LvCAё]VJs�\V�\�8@jқ���F��8��l��+S��(�h	�K�g����#������I�;�8��g����g��!*�%�2 4p�_�q���K6�X7[zW��=�$pj����g7��G�5���h٣y4*� HE�(Z��I�N|8�z�����0����yv���~��d�"�R��UpH�-�f=��!7�ۣN16(���ɨ��H&�FR�Y��>;�
�h��D�<5���ѳ�|��P�1�r�)���+�O{5�y�z�l u��L*���ݒe^�q������<���JAy�?�ה�g�Aj��u�r�R6Hp�_e��'h���A3J3J�9�����Xtn�H�q�U�]XɿJ���y��z�f��'n�K�ix�X�p9h6���L��)�|>RƤKو|S�E�s�d��3:v�4-��H��tiCu���, 4㯘U�q7T}ŵ\�1��,\�ϿU�U
�-B���Lm�`�؊����eR.H�[.F��n�{�y�0+�3��4i��A���w��ܛ|��S���K�h�;�s��*r������,�X��*�^;��
̕q�!v���|!\"-��`=G�dbyP/��J� ��,*�������(^D��r^}�i�G3'`�aM~�'�<�Q��s�����s�{��B���S�w~3n�ǀ�L��rȴ[�]ʘ���/�1�G��8�"e���]ʳ�޻_�D��p|�?�:�[�[/�㧕�a�M���ypY.'yL��=��t�j�X�7z!��QO�*z���������ā�/��"��)�*��U6���h
~_�on�X�7��x�l]����A�8D�ju��p�N���K��i�0�:���ޚFg�Ij������(f]�<���$P����a&�0�`�>p��]�}7�͙������2�2@}}��S�+G Sj�3V�)��e:P����A?m�hCS��N����l����`��ax���ľ����_������qQ��q�X�_Q3�;X\m���!�:����0�	XGPa�֩K���mB���`|gnQ=��9g/ۗ~�	MS �ؒ�V69�צ�}��Y���s�T0�Ȥ�E�BrN'�����I���xb���6�Qz��Y�L_�݃�蘽_�g���^�hi[Uo-T���3繸�t�~6�I,���-�.�t����K=�����.�Q�:E_�1��3��N���0����,awR�~a= ��&�^5����]G"��s�B�������!A�*����kOI��c(߿���C��i@=���p"mۻbY�|��X˙Ԃ�c�U��z��^"g��,�krZ��N�?	��=&Ǟ��b='���1��Y�:"�����e��x���(ҷ�Ӂ�0��� ��$*J4��o0�K����lw�NqZ`vد��$X�%[�@$������sC���&t.G،�����oS׺��7��D-&�e���3�r}��s �{쬏���lenB?!��z~�q�G�w��Ti'}����e�Xe�SP����3{a���Z�K�r|��!څ�S\��Y^����)`� ��U��������̃������"�>x��&�6G�Ak����u��{������6�R�d$d��o��Y��=�or����{�7f#y��ˀ~�S���|)s�aa�Ym0D6����lF$�ޡ��i��j�Z6p)?�(���PP1�e޶/�D�uk���'Jq�S���H�I���Y�}5"&]k��+ҿ|�����b�uB@� 0�*��EB�JX,ϒHgy�DA$���r�0��rxȿ�N���?H�6�4���nr�˥��L�͗ϰ����#��A���tܴ@5}7�x�a�CH?(�"M������ʂ����YQ���|���0~bQ��\���x�5Ux\ԙΕN�r1�7ju���W��� (J�v梼A�gz*�2�|nְ��WZ�0��M?��:I5��R'}���FjL�x�Q��*9���t�Q��zk�#�1�yt1&t�m�%�2t��#���f��ܜ�"�${?̾���I��\��(x���mz0�$r
f��.+�o"�Ƈ�Y�i���<�;'���,O���>��{x�	5�*C�P�p$|�:� ��� ԩ�O��@�Q�LJ���R������X=[P'H`�2�O��`x���(^@C �w�R|[�8`��d|�F���ߓ�SOa�5���>q�d�;�����Z�,KQ[ �$R������Oj��<j���~��p�I����<W�'zRn�0�U]2Z��`���C�~D�2��0(\ԉ7��'�<nܜ6Y���Ƚ��d|�bݧ�49N*��sk����Z�����⺂���ٽ;xly�`|��b���-H�iACŴ�����#X��JPp2�xv�R6��s��亯����jZɍq��/��j�\��<�-Gk#I(oKA��-�X>�05g��å׎�kYUQH�f�MP����[lM�����L�U��sTܬ��Z����_\�I������FU,���B" �[������z.��*��m���> 6cb萶��&�|Cѷ	�͛���|
�/Y���NE�<��i4���������˯��V�$�ǀ��}�>�м��0����@��ڜ��L����R>E��Z{�y��RW�����PF�=i�E7��v����`�l��D��R�j*���:AY�,��cz�Ø�ԍPl����[�o�nu�=L ��˹��T'����g�;���O#E�K4�wtj��a���	�а^lsg�sw��S�s��R�^�V��F%y����w.�c��5h�G���>J9swr��&z�O��X�����#�$3V�?`��ၖD��!�~)��~6H^�j#b�ɼn<�¬���y�DX' L��D-��Ey�"�ʜ��j��do�=��!�f�if3_�8q��J�At���rZ�A>�Xd�񚁋1���.~ڛנ�`�=�{1v9�����/�e��Q-]l���ζI������"�N��H{���T��~!�{�T�lU��h��0���T�;�X�#,]auk�[�Ԍ� ��k��1�>,p~��ٱI{���A\ש����'��䐅���BV�Cz� ����^#��l��oJ�����MO2H�a�V�Rz6����b�/{}+�[�j�,И&���z�Qx#B]�n�g���N�ZVyJYk(������?]���zgJ�|C����G^�M�a�&���%p���������K�(y6Ɩ���.SN]V2�@��3�4�g<;,-Oܞ�Z~�ԂYB��b3�f{���m�S�����H2؇*��kƠ��6��v�^x�~oC]�.?/��	�#��9zq'�F�#Ӛ���@ە�-�c�F��`,����jI�M���FO
$-��$З�zp8�^��9
ґ�(�ˢ�VL��F�{�)��ς�tn����n�x1L���4�(����7����$�]`ɍ�Ikn9e	;�_�5ob��gV�-l���N����-U_��i�Y��~W�W��������ł�LZgg&Xr��z����4�$�3��)��L9Ԝ5dg ���/�w p�9k�V���\HÜA�#��=9�2F��^����pMݧ��c3�+��d�tIg?�x't��J�``�;[��R�5VX�g{��I���D�.�㈝� ��M*mM����*ak-���{�tϡ�-]��/T���ީ�Ù����%�X|Gە�CI,mT\k��@�\F���o2"(2&gb�ǜ��.�������!k�oeƟ55t���孱#��T���c?ƿ�8��;�����BR+d}���;�1;�@jqk�H�_Sqh�uU1I�`�U�:&S,����8^��錣��ΰ?�����'�`6�Jh���w0�h����%fp�lU/��	�'Cr��i����[�OᭀfpKQQ�,>�JkT��>�`�A�o��s�8M���Χ	���|R�s�_z���Bxq[Ԍ2��[��Bb]O��e	l���tr4S�J��Lj�Ul)��؟��mh�W]ѧm\�A"E�5���a�
!����̐Q�R��ޜ-9ي��ʪ?�S�u>��u�ԣ�� )Tr�M2@EG`��_��އ]�{�a�;UIm���wE�m�v��B5F�B�;|̪]��lk��ǧڲ������o�`�c���K����R�M�4Ng=Qެ�����2$���T���g�\�@��)Ʀ�@�A*"
=���-z����a?����w�)O:)�	�x���w8�$Va�:z���E���
������/�����D�pqŕ�v��#���hvc�ȁ�|�+������'u|�>����=g�Q"|>���W�TBqF���AP�u�"	���UO46������%�cO.L�(O�D�M��,]4�ug|��Y=�ԔT$&��0���dd���`����_�{�������^�f�l�/r��]���Q�������
R�Θ<#��2:	���������ٹ��ew7�܈��+�r�X�\�����N�/��@�Zc��d�4t����rj����w5�&II�*�bte<����;��8Џ��%�����E��ᖻ`�>۬ǋĊ�#Ŷ�r�ᕷ�LE¶���� {�S�}����LW�
^�*5�A���ПJ	̦��G���w�Y�[S�_<N����������3��A�mP=n��\e�5���i8��ɡ��2U�Gx|~�л�/�M��$��;���C.���A�QU��Z��5�,���E�kx|����z�x�bl	�%��ͺ72�Vab����6���fx�k�om��2g[���9aU��n��㑂�V�((s�a������̘�J�|$�(xQ�U��,L{,� ���̙&�I�d�H�Y,H��#�\�Z�+K�Ϣ��:��y��X��"�c�X2����I�]el�vG��̟E�v���O9ǳ�+�FT�{�a�U�Q��m�ˤ���^˵i˼�:.�QP���,EO��p*p��� \.�o)����҇ژ�o��
Y ^��M����l, ?T��Q<ǏN*m߽"��V$^B�x}�p���i^��`j�,ItL�A�e|"��z3��k�ݼ���&zu�
e�V��);�)��(��j�� �v��B��@3hڟ�)s	+%�f�2ΰ��/y �EfUv����2��5���K31������A+�&nv���4k��\��4�`d�k�?�K&�l5u�1�9��0����G��Es:\��JC����Ê��lD:l)�����q�mcL��~_n�J��	��6읟F5$�N
`B�1u���&����H9/eDb�e[�4�;�"Þw_�'�P@��=���	�gRQ�h��+5FH����1�k���"����8O !!h�!��'����ˬì�Ϛ�:$��;~C�\���oF�Y������H����L� �֥�b?�t��s�;�R�������3Y4i�2��Ң`sՃ��Y�mJGQq9��*��(�������[&PM��T���uϳD�"�����.�����������5K�+�HU�b᲌�Y�Q~��R��$2^�U%���sg���Kw)�p<�(�3�e��6�nêЅbWEmd�c�5��l�[�-�v��v�����f�!AGNMDuX����ϴ	���߫��l��Cs}��uF���s��H߫�а2K��ނ��ܚ+`1p��q�.S��rA�N�`G����#n� �0��yQ/��H��$�؜�Z�>(8�P�R�����$坙ő=�#Y��T�+`��G%	�t��p��T1D��PN[-%OWD�G ���S�����?��6?��-��;����fH�3�[}���G���e�p-��'+����Vd�&��\���#:2*�]�^(<OEo�g_��j@����}Q� Y"��:g����f���'��N[HH�7WW��?�*X_^y�/M'��J+�v6`+����� ��1��������l��7��E�<P��)��5M�_~6�d�&MvLa/2�9	?]�t�â��.K�F��ٖ�7m�gL��O�#�՗���tC��ku�m6M%iec�D6��ƣ�m��V���ǥ�S{` K������~�%��%���I���DPy����3���n�JN��ݑl�+����*�H���P��
ʳ\�0 u$���23~*7X�̿��{�����A�6��AtÐ��BvS'���5a�;jv��ul�з�z����E��,�+d���NS Z!w��q���+�����
B��.�D�q��4��:�֔]j
����bP�l`�R�x~�æ��" +��S�iE���^o�{W�W��%Hs(;L7�s����6zU�u�ƪCYb�ď�3���� 4м&�4_H�^��^��X�!ȝ,�K����)��&��M��q�}�浪i��9p?�a�r �Uq�*��*���S�|eĥFvs�)��Ř�G�$��y�Td�	⦹Z8��tۺܳD�[�����")a Pώ�T%�GW*��GU���Ռ5�̥��JwW�]����w{D�&	�Ҵ�b����V+׼��I?��T��V�6w��6J�<�|��T��w�?���s��q�����H]�ǥu���AS�W.F1d��3�:��O�~�����ٸ��{�m˫�4���M��Rz�;/�gP%v���\��.4O|g �Vܷh;$���R��lr�nП`)��Q��F9���'�o���.v`!Vخ�F�MsX�Vу�H`-�6]/mǢ�b�# �)�>a�6ݲ�a�1���GMi����n�l��z�v��8H�T?�sgP�|��:�<%7ͺ
�}Q)_l+8�[r��a��	2l�ut�����
��k;(���("�{���엺��֋X���ZKm*�1�
@�ג ����;�$?X��$ED9I$S%B�v�,U��&�k"�=����9�\�����N�C@�3��nk�t��"�$��w��3��f#��i4L'4 uO,eW}c�V^�幓UF��HM��؛d��=���APw��ج��)��r����o�ue:��6��P����8K��.Z��d����q3>Ĝ��S�G���rrp�oJ|����t��Ǔ��q3�.
ph��(�J�(�)r۟5s���|�i��"�v#E����-W8��3(�T��������
W��%�BB�H}pzV�SO){!"�BV}���J������C���-w���Ad�}��7l�ɊO�`���T墻�IO�]_�1M1!*��Y���z7?����3VA�B� ���⯪�����q �\���;���+�b�O��@
�����k��p�t�YO=�����s�Ǖ˩[�.@#��9��\����G�vɡ7�kkN�u]��Q�k7X�
����/a���*�8Ƣ��Ty�=hO��D�#�9�!���.�L	MFuvɍD�����F6�Et%;���FO�ڥ@h���ELw�u�{ơ���I���Wd��[9W����4��2�� �=�x!�זO)f��/�>k�s;�n����s�xJ[��M�>h�&r%�9� Z��<����;K2�0�(b���"��������o?�t��OY̾�ڏ�'�����x��������$��t��^��6k���z��d�#(,�+H	oIJb�`U$Z� ����p�A�;��骹R-�	cD۳�@2�T���\a�@��PT�t�2[�c�+�I�Y�hyJ_7g��R�h4y��07Y �(`O�V��R�<8���d\���FI�{�ѳ����w���s�a)��
9*�eO2<�=�0�`#���#~=U���gka��z����p���l&,��d�]�:!�/�����P�>	��S�D�i����F�W��]���"����TFK�O	�-�� (�zMs|���d����J,��,�vw��<v�g.ro+�G+H�j0��L�1S�u�
�H�����{�+�&ӊ6��/�f->�>C��wc�����y/ΦFk�]��D^˗�&$��׏d����K�J@k�U����j��][3�4q6�\p������o�2R߿N�$��c��|�f-�kW[��	v�u� :���z}4�ٟx�%��5�w���'"@FJ�dvU�U#��+�&�.I�&i�е�5�Q��������s.�����它#-��SZ��]�R�ȍ�T��&s.j�C�7��C�G��I��&�X��x�6Ӻ��>����3�v5�Ӹey��Ӆ��a�e=���M���O59_���5��$>�-!�k�s���c��5�/�Kx s9��?��Qhb}��'����"�V�
��m!��ٳ<������{�CW���Kb|0+�5�ť!OM��9��X��S����#E��p��䔦Q?�)�&�cd����-�:�\������+�\�T"���H/��wA�葵�YA�J����Q��|��d�/��lh���� UEm��O�q��A?;y�A��F˵낊<z���O�/�:�q$esr�-��+7����6���\ˌ�R��2�x_�s���K^��$S���j܇���;� ,M�E��9���ĺx�b�ZBg�InAL K2OJ>�0u�Xe���|'�ⷛ��a�$*G��~���R�uZ�k8��f03!{"��#���x6<H]�ǯ�v'�G��r#js��4t��\�,�=�J��?��*�*�B����j����WٰD���ځ�~�	B�eK�p0]y�1�\2T*T}c�ʤ]��ʐ ٚ�F1��\�tn���6ʣa���n�%U���-�E�.q�D5�\��Je���ܕ��m����j]��_W�lj^?,얅==/�}.g���]|��s�N���7�T���HH������՝��w'z�d$��7����,[���+jVZ��h�nJ��z�8K�6��_e��>bC�i����PMlMk)K�Xx��F�fO�Q+�AE��-���j�v3��խD��D�u�� չ���l����EPKS�����D[[F�H�N��Rs_�ɥ��8�ܻ@���y��fPuE-���m^ �ᥴ�C($=Ya׍�:x���%[Eu��B0�W�����
D��6�I-Wr2�C� G௻7?�j%�[�D&o�밙Ds�:֊���6�.A�/7�c��.L^5�]m_�`Ã���{���G��P���V��j�qMp�?x�]��&M���A�"=�P�R�1F�h�s�@����Uz⺣�V<�&n�x�$�AT�/N�d��"{�4�1ΰ	�6l&-���I����L�I���ǚ�#(X�x�"J�N��}#����+�Rjb�p9�fyFO��$__����m�4U�]�1B �ڟ�l�ב$�Jk�0Xlù(QW��m���d.�?.e�/�6m����$�F�D��F�g����oȀeE����y#��!�+�:}���vk��":��l&V���j\����ۜL��o�#ֆ|i��;��C�UIR ^�k-_�T�}ec�R�bH�-�_=��a�`(l@	6�7~T�(D��4N��r�T'�U�G��f�}�o�t���A�Jh���2b��|
Wk�W�V�������+e���� �V���[ı�#'��k��oL�hn4t�ئ��'lS��w�Q���΀�r����$$�;3U�X5�Q���i� �L+n�GU�]��SvA M�58��gm4�l!��/�$����a���Eb�\�
}���;�=V�e���Y�I(W|����~�ަ�j��A����7�_�BxFڨ�bV�=���p�34�Ǖ�=h;��j�:˧�$/l �QD"V�:c�J�v+<|�G۷�4�>��Kl�2(���![����V���_9�M�qE&�-:����.z�&%���Iú`&!-:�?���A7ֈ���eT��l{d��uhW�� �8��` ��� �+��;�a�����T~s���fA��s�b��QV3���u�q�BY�	 M��(��$Ў�u�y�TJ�g���SY����PU��]Ch�\r�@ѫ�m�6)��ZTn��T̙��b�\�C��W	37�ӣ�̷;HZ��(.(���
������EPc��@C��Bp^��M�D�,���������X}�wM�&Mh<�َaN^�r�f� �1)��F. nHȱf��$Ow����Y��ʅՑ̚�ȨR��f�"O~������E��q��Z�����{�cU>�rU�������V��hB���8��۩�l������ں~�<��Fg)TR.�a
H	Hu2��3#�g�O���P�RJ${��:b�
s���Jc<��"f�� G�!��5/u�߯�����b�m�jT����3R�Y�!�����(�&S{�#���]�$��L1���~ I!^�B�LPޒbm��6s��!Ì#*�f\G��5&��PR2ɫc>w;"�h��11��+[eѮ,]����
�=z�4H�QC�4�d�H�����v���R�F&���Z�X��ˤ
ۇ��et�.��N�8�@��i}��2��r�3fG6���.,|.��V�v�$��<p#A���� �+��#OT�L��������ܖ[q�|oc��f�91
�±�@l���;k컱i���]��Y���o���_�!R�����,�j�B=�n��Q�|Gi|A��f�T*@�X#�șC3g�3���rk*1n�CA+6#�=ZP��qTf+�Eއ]	�$H�GW�D�K7�t��g�S�m��JwL)�l1=( ,'o�i��lGh�gS3h�b�ef��ʣhq���+�*��2��:��R0o�W�1lG6K��E��yo����-�A�[���F�l'>�`gs��Q7�=�B�	Z�`�YȒ#�y8�d(co��+��p���$�>ـ6q�4�w0~��,�u�g����c>��#G��Q��f���)��;sVk����ɞj�N�L��7q�E��J~u�J��E1�Uq��,D6��
�kϵ>�8e���r�A�&:�����%'��"�D�������ۯ���c�;��a�����e��sna2\O9^&�a X�3R�[�jL��)y�e�ŰH�<]ւ�Nx$��py1҉�/չ���.��v�"�O����pZJ��hZG���=�;I�1���l�+��5��_�^�]�/M�ۥ^"r�՚.�9�����hM�<R�D�K���/6����� ��{o�OmWz�����k��ٸ�P#.1�(��3�I/��U�H* ���{,�D�%Z��[y�M�^�KWh�2U.+�3���#�����v�`�����%��#�x�bd���>�'�V�1n�Ƀ=����\x�<"o�R��V)J��o��'��k��k!��� ��8�X�ʪ8�g5�\=2���Ű>S��ٙ�}�^0 �Pe���MW�x"�M%A��:��e�Kp�h�&�G���08������w���f���]1�B\p��!i�#�EW��l6�s>�i"�\��{=5Z]B��9�v�l�iL�NA�>2M�G8fΗ�8k1�G׽�C$�u�����-�8�\A�#L���-�z~^����g�z6E�<�"���h���]���8"��PU��l��w�)���ze��+Z����f�$���'��Z|�uTNgSRC�����s�h��Dg7�d��������@4���W �f[�/?��䉡]�:[�]鴯�#WS�?�%�!50���>��O�Lػ-�Q�#���^o�X���m�'�.(x�	� r�s��5��i���T�g7hW���'���<��ً�f�yV�-U�dmrӀ����Tm���D*G�]�u;�@�绶[��v�>F�����W�����nt*�ʦ�<߉�1��Q`�޸2�"9V����7�X��+���T>�W��I���A�*��w�� �Y�M�K�)$}��<������ݨAP�)��C��C�����"ngo%��~4�Pw�S�_�vf03828^����sB�Jγ�|"zoMajvV3A�%@�_=Tt�66@A]�T8��_G��d���@{����=���r��}}��(aq"��ĝB�ge����Y����<�&|�'��tQ|��S�%*�b��{ ��#3Nֈ�J�'�Nn�o�.F6���d.���E���I���a��(a:���*<�\��?i��	M��'��S���cJ�LFs���O%`�0Kg[J.�dQGŃ��.����=3|�+�"�S��bl�県�G������p��� ���u�d��cC��U�h��vۣ����7 ��!�uS�{��[�f���'���ɝ)�<������®El�\k���L�[d�'��-�����s$�V�jt�49m���'����!t0��z6ڑ��|V��;�&�>��H���tR��-��f����]��&^�液���Wc�{F7�z�v���4v3	�=���Jm����)��G�YJ�IԹ�?Ig9���̬��3k��F�T�p��zN���*�[G�&w��uF���YP�ř�Ѐ�7X�����]!Z�H+\�ף�c�u_LK(x���J6�u���_LQ�%U\�e�8�M�|�2Sʢ6���]���-�@��Ƨ��ÄKz�e�٭H�( �-�o���� o��h4��mRX�J�ǈ"�r-�O\[�`Rh���t�l7m�`KTgWNE��&�����F�-r����T���6�a$�����d��bS.�n'�eA���j�oMqk�w	&���g����+��M�KtP�4}Z�A�Hޏ���w�Ϸ�g~b��;r�Y;�t2����(���o2�~)�|s	��֒Sh�}S�]*	��d�Vy^���*!g��(��4�
�e9!�)������}�ͷ�*�,�s�{�I�XH@pj����QΥI�����E��,�����M����!�4F�ϛ��9<����iJZq��?�� b/ ���#���Y��)3.��R	�F.�)��/�&) ��L�*qA܏�Z^U��v����{��]����~1a~�X����\5VK�y�ժ%�)��t�{u�T�Ǐ����h��Di�>���Cm�!�O^��58'�#���JSz:@�o���o���p���M5�A .���$��4��'�3J��OŁkv(���R�^��J�7	�ى����0���OV&���hT��:O�'6P��G�� �����ZF	4��5d��~�����s���_m#�<�JJ}{��+W�D��#��k�B� ��[&CG9S}�4������Pb��NK\3.wU�O}��tb�k�}n���bX׮Q�G�Tc�n�Yʅ���q��=������;L�6��:�b�0�Y���b;^���N��a�Q��*�-6���'�������� ��~���G�xB�������ώ��r�˸��cjft�ҹ�e�ex�n��܁�˽����(�uП-X^D��;<?#�Ź�J�0�4߰���pz�AAi_\�0�̎ ��Z�T9CIt��߇��'�|�=���}�O>�
b�(p4Jm��\�n'��^�D+
��8�=�}|�Ύ�$��Ջ�΃ԡ�;���5!k��L��m��E�܃�v�B	��b8�]-��@�a 2ˮ{�؎t�0Y@���_� ٠XƳ�4�s�0���=�MI~�[�?� ��HUu���`J읾$*�#�=�;���v˭�[�b�r\���� �� ����Azm}�b�����@N�y/�L^LQbH����<�k� �c1���������kX�1C� �skd�*}F��q�}��4�}*�B�nI|��&I߯��/��*��^��O ��`���T�a*��?���&��á#�Br!������]��</��P�4�$�W��$�mPb��N��o/<[yٜ?!7*,���<x�5�/"�N&���4�� �SR� L��'E����g�|eDP��*�Rd���/!�H�*#V ��Η$�1͝n/��Z9��h��ڲ�u����%E�@|�$q�t%/!�5G�����lA�wp^\ZAG��x�۲��Hk��*��JS�f�&Z.,����P�ӥ�K����0��Pn���g�mUmSe> �6s/=_���.�����5��sSHY������*�ʂ�m�嵙玻 ���ڜRgc��^����u2{|������D6F����a���^�}[��-�`r�u޳>iu1�(��Ar����鍛�=��Z�I�y����Nzʗz�lk��Ԏ�{B�BMOj�nB�ƀB���{��dBDf�x�����20�����A&�Yo��;�"ns����yT�Dd��q�Cy4d�@��r*�nwT~޳R!���z��Gck&Ou��QC��K" 8��5\���-��Mnzk=��7�	~w�EJ꿼�$��3�0��7a���G�Sw����1K/��4z��v�z�xjע���3�_���Լ���5�)�4I�
�F.�̒�֠�@���*\?\����4�	,���B�_��X6j���n��F�/�Ln���q!Zˮ:ݡN/U���4���kb��@���]fwgȾ��w�rj�V�?�����X��A>��Km���
_7�V�EF[�Ox���$���n��{��X�H��,v)w�!I����%ã�I=���LfpP����D(f�=��C��sj󳋘R�Y�-�J��� (8�l=hI�L�U	܆�(�J�M���ְ�M�#��}��(�VS�j���q��9n8���n��^lq���awzQ+�~!f����#�/��3��ծ^�+P����3M���S6�7��P�'��m���f�"r�&�
J�}W"�R�j�]��;���i� "bD�+��
� �yD�F�[c�bN�	H>�	�nh��DA����)x���_��j�Ĳ;����8��?nKdVY��{���/��9�F�!=:�0[{S10A�cE� &o*���&wċT0�l⇖5Jk�#ӨĂ���,U���b7��)��J���~�ި���r�3hjV��m0;��^��	�fwQoSW���H8�&�����,�� ͭS�F���Ѩ�ϟ�sR:�o�Q$�I��XM��`��.B]���嚂'|���y�%h�uЧ7b���B��飩?b@�!�X|��+��4�W���&�܂a9�J�z���F�9cb��1��T��}�L���ᗒ�@�L9R�CI&��Ly�6�S�aw���^�e�؜��ғ/���j�,1,7��y���jA-�r�UQR�ݯ�8���/���E�*'����A��L�V*��%ʫEw���=����W$*j���.-�;���dZ�"g<;8�*�;�����x̎	�s@ˡ�|q� G���+^�Вr��~�Y���=X�$$����,~�h=�L�ϒ6i�Ǹ����;�����6w�\���k�S,w.����j�����fT����������u�'��ӕ���%�BN��ľ�>N���f�����ẜ������V��4s�|�v��FL��|��,	���\"�?dn��Jx;�c��U�fmk�=�h@�+co7�ǽ�t��G��q�r�rw�`�|p��X
��L'�_ϢĈ{T��?]���o�b�J����wr�\ߘ�V��ث#Uv1���������o��ھ$<x��Glv(a�t��ǎ��P��� Zw�6rD�$�X�Jߛ���V���F!�/���`��ʨcK����A�SN#�?��oǲu�L9q*^��B���M����+����<_�ܦL8�p衇��HQ�E��n7�+��F-Eve�+W������\���x����=�;\E��Z���rn>�I�Am�C�Wg����K4'���h^�3z׼�����	4���zR,F�/�cFN�����IƱ��N��v*������������P*$+J�ET��wl��J��7H�/>4'ULj>N.?S��q�^����+~]� �
�C�vI>Hǖ����Υ+]�ډ�>�`�!�	���j�ە�wZ�I�gL�%����Aݷ���3Ƀ3̦2]ﱙi@������G���4��@.��Y
��>�̻�3pk%%m��~K��n��O�.��$���I�H��R�#�RcR�>�������������}h';�I������eG6���'k#�sD�/�"�c�k?�Z4���4���	���-��s�DX�x�²�Fo�:�A�(��+��Pa�4O�7����`�S�o�.��r]^qNc[a������}�a�i��S$�J}�ŤO�\[�CZ�g��jr}Y\�S&�)�/[k]����G4��W�Eӎ�v���)NF -H�A���ژ	��y������Ġ�:H?م�(-M�1r��kC��$#�̆Ƶ�ٔ%��ݼ`��1. �S��i��Y�&a;R[�?P0'��9�S�Mf�����94 �;}%��'K����©'�N��[��1�l�z����y)�U�"�Y1����9M����|�ޯ -��V{m���S�B�������֗?N���g�-)�1h�k�ߘ@	����g���4O%Dt�n���Y0^zZ�C^Tޞ܍gc��Z]�cbô:$\`X o���ל�0�O�4�w�MKn����$ˆ{��� ?F��k��7��\��Z����C�e�1
��C��}d�>�{�K��5�7T6�:B��~~~n�1���-'����on��hJ:��	8��}2�!�Y�z275�6=�Đʩ#�We��*�M$��f:�ϣ ��4֚��&(���l����JӑL`����T����.y�ۋ�X������>]<��%R�g��\��a��ΰ.jHq݌�t�7c�/�/$���c:�`�v�s�B[�t�kh��1�
������[~S}ݔ�I��ݨ�[��5-�y2*��B��?ނ��ƚ��cd���5��;�eC���Ns��Fq;�S��T�����B�6P�'�=X0�a���=٭�iZ(�l�p!1=ǝ3�ط1]�&��	VM!�$��x���0�⒱���vN�f����(|hu8��F��r|� ��j0��^���w1&P5v��(}v��=m���<'���,ƂK�(�u|����L�<!� :8�F��{��Bl�*(�8�bяs���d�L�����<�8��:K~�]���*��K尩��2���y8�����������*�����f�]�N/ze�Z��K�J�g�7^K��>�*]��v��,x�8lӍq�n6I�kbG�TR�{��M[�>�����uY��4J����e]�؛�
��d9>%B\����uV��w���7�R�W��Ƨ���#�lt{,R�d^BjT������Z.n>|����� #��ˣsZ�O����v#���qPk�H��]�W�U]ߐ<��[~��ͧ��ś�L�:z<T����@G$+A�Ib|�g��P��lQ���������*�j'T�����~ ��
�nt��\�����^N��Ȭ&
�B����k)t�&b����=�4DI��3fj��MVґsX­x%XpB6g��(�A\g%lėУ�_LՌ{�<w����d��gm���;�=����@�Ti�����T lYs��}&�6u7EE�gks��ce�i"���Y=�z�&�- d��rS���y,Q� să���p኉���~ng��N��U-u`=��F ��C���W��ͺa�SX������v���ۨY�I�J���8{SI�8�[�%��E>���OD��3�K�� .;We(�"���y�eHXoh��U2�S���3fPs�Q�h!��|I�N�k���w�U��EA��Lm��U	އ��6_��h�r�ϊ�.|;p�|k����L��^y����^�t�.�n��Q�pՙ��h���)�W�t��/bd
��q,\�m�G3?V��I�s���\&~����;_����g3�C�,8>��̖2��~tGk���]������Fm��N-�y��d9J�'�g�~ކb,y�*�;�~�������w0]B�o�&c��
]ܼ]=�C��l���nɪ�a����LL��ex2����k�;�����6����4]2ZZ��ل���Ǻ�AL��1��V���x�A�>FW�-L{�@�d�'JG<�ӊj���ȊV �z�ǔ�˜�P���הX�R��+�\qQ���� �f�Zw8Ć�t��_=;A\����r!j@�d�0a���Mӂ��g��7d��&�J X\�{�x��XGm�����<����SyJ��"BP���PԱ�s�Ms=,p�kb�ZO}���F���S��_}I�;����u��f4��J�g���&r�TG�!���W�B��EC+6	�˒��ơM�(�K�o2K���Y�Z6� ��㝟��
��$��1�ϾHT���~T1f�j7�?�	9��y��9}�w���qZG�3���!�r;`g��@��8u�P'��y0k�4�%@�����>э�
���T������}��6K�ޗ����\����@5Mf�D��K�b�82,<,������yҹ�㲷5NGS�l�^ѩ�"�0�Њ�?>���f��V��4��-ͱ�K��d}�ί�v��e�w%qp�u�
��.׉��-��L ���bm�7��1�Rď�'�^!�%��{����?�UPd�h�-@U��h�ɜFo�D��N� �PU����|}�(IW]�Չ�����L�K#uFvg��n��_���I-I��]��#�J�4a	PO�ͩRA��gZ�@��T�~�&��{�!�6�vp˓x|��1�Q�"�|�>W0��W1Lz���qG=�&�d���J�T�H�?��&����\θ��g���
$��ϒ~�W1h�0�ޡ8*"������s�a�&�O9������x�eN�jT�9�|=̷@�ޱ�r1X�9�A44�X���S�^�%$��\߽�*rs4Q��R�{�̦G`��W�^�&/Pt��]��(�IBP�
�"2 N��^���:�
C��>�>x�֊ZY�Ny�`�V��ÝV� g���+��6�fR����<��t��0��Ȳ�ߒ}㾀:�9yW���I>��p�"��Zd������/��&�"* Ua[D͎��w�	�锲��~���sjMΩŹJP����M���8��Mb pp}݌9�@�[OE���_���fE���M�-iz�Y��2���AK6��h �� -��cT�"�]U���� -D;�ZI�_x}�����j(T1	A�=|����[�'S믦�����K֤��i����W�qĮglN>��k�wmK.�Ԋ�aK^�v�CO��-L����˹]��l����Cl!(`������87k���~���~��(��yA��	���OnS�V��5��U�t _BU1c(� V[Ub�63�|!-M�� tK'{�[�-�ƭeܵb;S�3&ÿTAP��4BP(�\b2���U}E��JΉD���^��� ��8!*�������U>�s��  SFmlDp�{\�C�x��\^�H8�n�p�	9�<�p�Cɒ�8�U�[�\�Onˣ�ءI��\tk.d��V ��j���<L�Cx��/�:+��q�,��X�J	Ȟ�]�b�(a��GXd�U�[0��GU`xMCN{��-w��/�[��]+8_����(q�Q T8�����9�5�v����	�Y���$O���o�V��M�+�:/z*�1F�Q8�rOA|yVe�	���Co_���t��M�߂ͨ�Ȕ:W7�PY^�o���gz��?������'4s�XS�;����!b\J�Э3�j�`�ɹr��ᖤtr��χ��㫧-,0�<)I׿��S��J�m�'t��P	�eh9��=��J���8�P6<%M7eJZ�H������h��w�s��u�ƨa���S`�x,�Eo.z'$�ҋ����(f���_�`};�%	�U�u-G��\FP��GxX�X��R�����R��&
1 �7,�]b]�3��/2Y�4劂���Z��P�*U�N]Ss�;t���A6�"�~,�wV>��|���^w�|~<���C�j0�8�
"yf Z[|Y�^ыw�u��h���������3
��0�<�c�q���q�\�5u3Cf�����y���-ꗻ���"r����0���w[p�ִ�e��<BEӢ#i�\�ꑝws:�|���eW�:&�����E؈D"�L�&r�i+v,S�F��b���Eco|�!����va0���c��	�7�)�6vZ�7>#�ז��ڱ�@~�1�P���ÖQ�>�"�*.�f�jJ6T��-ڨ�����9\K�-��D�N�Nt�s��\����Ֆ��.7�Ue��HY���pZ</���0ۏ�����r��G��JO�U�j=�p�Pa>8Qe�^޴7vB�	>EM_b������\7�H$D������ˠ��fS�ﳭ����B+�t� ��!1�ԭ�T��h{���ֺBL�/�HS��y�w��.W ܴQ��;G�;}С��9�t?0<69O��[���{@�[��+N'ښ�	~_o1=a-��"�~��(Aw��X�\!��|�2e�w�1y���) N�Uf�^`������e8�ĝ��=��:TN71a�W%|Ot����90�*Y/1���{�jP��O���w�l���b�jR���ɦAE��!��۴����wR� `8������P�Ԅ:������ѣ��2��ߺ�߶��2�%��1$4��[eÍ}J�p��k#}��n5��=�m:�H+q���7{%����虀a������s+���(e��w�E%�}����m�IVm�
VLN��%5X��rfdun�Ӄ��Gl��_2����٤�$k����	�j�����ah�i�k�&�q"5���n�A�q|��7ZI�TF���h��*��]�\�Ko�%9�%ɔ)'}˞	�gzȳocD�V�_�
��[���"9������I�T�+�:���4G٢tkV�)�t�����O�ޓ>�&�I����������lJC�7'S�/�G�$�ӀLH� :߁	���.��N-���nj���I�:G��)�gml���E�5�C�u�3��Ӯ}Nxu}H8�mI*� �ɴ��kr���q6�������_�����<��I��}���W{�ȶ��(��2��v�$�o����?Q֍W��=�ܹ_Y�"�5N�)����(�����x�Uୁ��M���|��P�Z��&���IW
n��^��S/Ng:�:+b��&�8���d��j��?����X���������Һ�eİ��7?g�����5a������΍X�Z�'���	őP�Ϟ��Xឨ����<���7�� �ϝ���S3�/��_��$Ɍ9�lg���i�#q���/<�hq�)��@A��i,l3��w�HC$ޘ�o&����x��H�ķբx[R������O�9�F�׵�L�c�y$]�I ��k�/q@K���¡����A��A�{)�yz��p�ƔJ��O̯�Tz�+���&��>;Yw�x��ߦWvܷ�@~�h�}V�C}oxf*�\��R(��z�t����G��p�Z�'�s!�8��/�=MŚ�R��:�J<� �M��������U)��T8�UtO�R�N�,�����%7��rɤ�ĥ�QW�!�"���'�#�w����^�O!,,X�����;�.�a�D��ǚ?4�<���Ϟ���V$I�(���u�]@��[�ҁ�am,�{1���>w���8��C�<.�?�zO��bYh�1zRv5 �S�V���f����#���߮��_o��"�A��$SsA4$<�s��m���/!d):6�1y/Lx�栱�f��s���Ng �{2�?��m�F�W	��[@&��~ge��p>���yiܼ'�-m�өZ�=2�W;�gj�� ��5��_]�^����x�����ߪ��!پ���85sc5�␋��4�!����LtzS��y<�	5@�d��$�%���M�;a/����ro���-%�2i['�b��y����j`Q����,�δ��6��S�2B�K���\"��;��!
d�.L1����6���(	�������� ��TB�UN��h�͉���ZĻ�����n�s�
HA���_���ʔ�x�8�������s	�p�0�W���2^ڢ{����׺<�W��e\=�7� U��1�\��<�T�+�����I�!�^d���#�߶2<�1���+�N�lL�
6��obȇi%\���$�huHl�E�9x�O��F
�AJjK!'9��a��ş�w�[Pm܈\��BD�Xl��.Î6`�!1c̰7�y�Bڰ�V�zX�B=zd ������_N@�"ޭ"
���C-��坌[k�CO�)��B����]*�A����F
@���	2Y�����k�=g��oH�e�u�.��}d���<�D0�̈́j�<P��r��,X@�F`�� �9y��t}��sjCnw���: �n�W����]!�O����wUoR�E�[	��8�Ӹ���xOt�g��IJd��3��ӣ<��s�Wb�
z΄INMj��;����"ӏf.^�9��Fl�Z�Z;U��b�o�5m=�C6�#I� H.>���D���jNA[��p�ZL�1v�Q��\�ѵ�&��!`A�V��*�Jt���~4>kH�bLY��Zl˜���hm���u_���tfSm�4�i֜\ġ /�lg)�lq�����V��K�͖�p�*�ׇp5��˕/��F���,�3��h����Dm���Ζ�~^�G�W�3
l"N-\B�鑫�|rs����وc���)��P�$x=���ѠY��ܦD��y�����zaAMh��s^�3#�h_��QL�����d��Hm�S�5��޹e~�r�|���3N���6:j�꣦��x����p�V�7H�]4 ������JN��bm%��3��6?����b$�5ͽ.QI��(�Z��359*q��{���B���h���JhAҰq�0'����̛��B�sߒ��g��r���e���MT�)p��
�L'����^�>��?E�p�)�fG�S��`'y���y����]�3�w�[��}�m�p*�@^۔�&U��U��*���Y�V$L���2o9n�4is|
��u��E��]��?{e�s����^!�4��쏤N;�t��,�[Q u]�U����������y�ta���XA�- _�7�g�;���+Mu�{g��ö�Ƥ��[8���m��[�}+�l�֛7G����HO��M>��t�>��9�g�}�O��L �C+Ϡ�9E�Q��
��v��rm� ʫ�x�h���k�S��)yܚ;��Ȝ@bS�J���������@�������BM(8��������e�/�1�h��`\#m�0Q^(��QA#��_��y\Ke@o��S}ŌH�u^�C��$����b�lؖk&yHE�1h�N^��K_�A�oo�V&q+��XX�Ƚ �S�/�⾱Ѵ9(��r8 +dZ*����t�s�a���շ��"�:�C�3�)e�JA��PI
X���4y��?��M�Joy�6��F�J�^��"�<�ZI� P�!����怗��G7�"mA�?���}����#��۩1Ĳa����>N�J"�jB~b���#�i��8�9IFiasS�����L)��RE6���8�!�7d��Q6d�!��:Ȕ��z1�#A��=�� vVi4�j~#����"�h�I�ݫ�z���bG{ Y�806z!����j}��~+�\��:~�GY�wV�/3��{����<�����]��=fE.<����8���t�����`C�;����e�S�(�i����SQ����#���U���r.���2$E�B�@d���zF���v�4N>�k�xqWK���DKN�o��h�|���%@T�a54z�4�Ϻ�GZ��;�;'ToF(�qs���W���D��.��9�S��?�3�PWϫe[���D�t�i�+3k�#q�pBԕcժ���.	���W�*� B�d�.��?0(k?�~�Cc�U�����������s���#�%����Zǹ�=(��F��o�n�L���܌%�il�
>��D
RRn?xCW��	��>Ҹ�˚���|�+�D����_�K$�����C�\�����8RA��չ�'�?���"�p���Y>j���Y��<:b�f|ʎ���+��5�1���n�x�b�0�/s�Zx}I�Ih��=S�6�"��3}F���`dl��	�X�њIx��ds}ρ��rlś?/A#%.:r<'��e��vl��e6y�w�4(�I][駑���r�hor�@���� �.��c��z^�n�Ra3`�����1��L� E���UI�s�~jr�`�T׫��ۇV RPU8Jke�)��J=��2��C��A���ɜ��N�w#�q�7���������fR�t�V4��B]U"j��`-����4��ڵ��K`x��/���*+��+����qۆ�[G�n��N{�?d��.�5(Sm�&��$�i�~�<����(�����#7�X2b��!�=9��T�1���3y��M�݆� ʬ�5=i�U�=c3���69{:t�,yT�H[k����w�V���b<���P�
�?�.��2-#�S��۲�.��č����I[t=�M7#�Υ`�$[j����(�pa��1D�*�~�,����8�	֙���1��J�ʺ�T�M�}�Sr���5�Ͽ�A�b����h���@� ��19`�)H>q����^�;�+�e
�,�N5)��fC�=|:�<��C[C�nP��ygF�����[t'ߝ3��"��P���4�Mp�{�	�i�#��|����a�б�[v�e\�Y��y��`VZ?+�\�Ox^�T��ăd����4ձp�_�Ҷ�t)6�r��^��o��?����15룙���J�\�z��#X���?�*kuf��(<>���V�p_�~�@�o��j�vq��m�� ���?k����+UvQ��k(x1P���?{z%�`dTr��`9v�G6� @�>��N��J1I{^��d��ƋqSt�Q�ى�#zG��6e����S�jF�=���V�7C��	�Y�����y{�%�ڎ����|���	�jI�&�1oI�9J0��(�i�\1�Y��OK$`�n6���.�uSsy��dU�M��S%�8NS겸�z��C����3L*�:���Ml\w%0�W��v29�i|�D (�����AyT�L���#iB��N�j�"��t|��	y���Ñ�T�ȴ���8���8���诶3��H����<�w<�i����\w8R�'=����"�ؒ� �TK��p��f�����P�>��"�>�\M[�XM��5����`7�(�Ýs�M�q�0S����ג`�T�l���切yl��Eg<!D
Gc��_2�h�ǀܳ͒)W3��ٷd-�*_�n7f���U����g*åc��o��J��!-$?IF��&��Y,W��F�	+)�~�b�%Y��͐��*�$�o��������n�[tń�7F|j���Pu���cL6���z���߇Mm����q�Ip�&�?~�@������F�t5]2~��n1�w�}����zc��*���4�} V��g��U�0��x��h��#. Pk� �������?���wD5H�8DB����sC���W3�L���tx�h1�/xy�*��k�S�)A��&��	�!�*��w<���C�U��G�.����?���G�� !i����J���u�p94Ц�K���BeIW���-%�!wݣ�ʅ>b1w�S9Fc��� ��+51<�A��|:t�
���{��`�B_����#��	b0T�%�y��n��W�E'>x�^C�G�V�]��q�-��g�c�����)��ďa�{�l�������j��ݕ�0�WG�M�k�E����˛�[�0�-��K?��������a�c�8%9�3���kb�e�2ͨ���U�!�,�<|����o�3��/|%ل���F�~�RZ��X
6EBp`�X�D���]�.�/DO�k�����9v��d��ź(sՠ�E�8U�݅��R�>*JV�y�A�?�	���.]�����P����&<DLVU�p,-7^�����7ʻ0�%.�O�ʈ��:����!�81h��.���O�v����y�������7g��:2���0 ��VR9���V�̈����  ҍ N�ä�'�a�8�s��M�k�e�C��d,�d�2��=C����>k�Ƌ~�i��1��S�LN
�`�'���L2VЅY0�I�&�����W��B:?���ɘ��a�<S��>=�����jә�-��t�������Ϥ�B���ۏ۷���j܈h����7�H���4�^�C�ؿ�=o%c�.ݳ�X����.�����8�i��~:�z<���r}C�Q�F��rK������OqBZ�"fe�B�]|y<���&�ePL���z���mE��=7�%i�|q�&�E��؁
�GN���h�.�g1�=)���n{��/!n�����T�������~Tu�K�ܕW������C�JAB���Y�J l���#��rД/E��~��@�2x7Oq��UjZۼ�~S�a�T`mQ����$����5K������=�!��]�~qL�>�������A��*���*�S���S��t(��rY��tOzp�ȫ�筢p�JxN��T�<����a���]a���U�E��!f1f^Ӡ|`Hq����{~U������h^!���0��
�i�����w�$m���MC�#t�nr�;�ҽ���6��`���f W.�Y*V�X��N�y9!�L6B�.�}ͫ�Q�/o�~�r�]ȧ��rK��_��{��Tz֤�����T�:�~9���LB�K�z]��q�W;ccD�@�v�~�cN�pǰ[jR�'r%���;���^�2@P�q+$��X�D�-���~���變��V3v���frPhb��'6��̢�&�]ctwԱr.���h��K����W��B+�E�e �]�}D�b���ؽ�ii�X"�Ry�"��W��z%��{��nqS���;�w�P�=��y{�]W&����y%�sʍ��M����8�G���R>�Z��`vG��Meύ��ĽE��/~"JG]$'[,:�>�PѨ��xw�'���RV��k��6��{��� �ޔ�OT�;��U���������Z|��6�V�Z�㣍�"P��=$z�N�^o��"u�g���c��r�%]xB3��Rg�E�A�I�9��G�A�C�W/0>�¥��f���C[���J�D疖"��@4��(�<Z[��6�1U ���H1�c�e֠\r$��{�8C`:�i��.m�X���*��zd����Q�&A�}�?a�&��!�N����l*�м�B�=�����`��Ƚ)v��K��*�ݨ$���;��~��gu&��
EҺ׺W0\��ɤ+��	B��(�f��A�w��Sr���t�У�K��yP��L�*aM���ܮ����$��M��� {3�����?l%��EA��˭���O���8���r}z;��(�x
����i�+���.ش��Qa�b�̓&s@�����cg��XNHfwm%	HW@��*�/LY.�ݛ�g���O�0T�Ʊ���k�Zŕ��f@�%�� !DH��J�&�/���ї$�.?������A�}�RF�k�w���M`��)|�]���~z[�ʽ&���GpB{������9;�;�x���3{eUȶ��fce%y���x�Ԭ��O�!��Z��`X�~�U��Hv]���"$p	(̔�������u��C#��@^�>����wkX�,��p��oЎ5�9���g��������wܽ� �n���`7�oܛ��Pgo"y�r.	�T�~�rY���?Z�\=_w�>C!���҈-��t��嚥69aD�>=���� ��izM?2�~�3��hH��M�5����k	�.YA�� �������S��Ok������dX�*�Je���s4����YN�{����G0�*��?���!�r�[#"�' ��hw�_����΍���I ���=�}Z��hC��C��ʷ{q�� =�T�y��J�eŧ?؛��8A��'q�g`4��lQ���
��2	��!��$TF�����$�����$U��&��C�f�ɲm�:�����R��H�l �8Ƒ�ZY3��I���Dd�Tzn� �Gp���AY-�o�abe�)+Q"�b�g]�U�=��*x|��c�:}D-�5���f�N���$bp���0T�Y2�uH�;I����8�r.};�bm�R;e]=�h�@@��K���L�� �ٶ�4��ƈ^#���'b�n~~��|l�R+��U"����EO��ƶC0v�_d۝�$L�O�<v�8��ց�*7�1�B�]d���=�h���Ʃ6��V�DdGѷ�j��(�h��X��-���.T��%�~�t���=���'t��(�"�%�f�����gMdg)zF��$c4��A'����m�앍���ӎ���
/��J�Nι��Rڀ�֕eH}p�h�J��޻ܜ�z��v��W񲧭��e���ǆ_H�0YO��XW���`�ɾMb��π~<��$�9��t*�2��9ۦ��>g(	a�g��7�o�aiY;�/�*'ȅI�3����Eo�j���gF���<nޥJBhחLtMB�փH �8�a8�+�&��c��.��H	�{Z`y�����\�"$6���f=�];W7������,c��(*|��
��$��Ә�2o�1�'�&�8����g�N�����gy�w�j�J��_(mUo�|��O>�H�Z)���4nf�
�t����׵���|�\)`W�6�<�Yo\�x�a�$M�ICF�](��ռ.y�K��O���w�f�ʤL<�3�>5�Ki�A���x^�%�zb*�83��byT�X�%����'��>�P7t�Pj ����ֈdB��5L��l���s9��~��K���[�	�r��.�=��&�A�.[6��;�� ~��>eTztj��g�IZ?���I?�	O{ENB�\5����Wg��̬y*����`=��Y��Y

�::O�Zv9�!����.�G����F�B�)"-�!�_�ɜI��V����݂���5p��}���*����%����T�GQ't)��Y����M�Η����p�f��<�ۻ�
����d�J�b�֔�O��:��`�XuS{�^V��Fd#�!%0�AH��Q�S��g�bY���[L�iZ�ɚ�Zш+��h-�������ng휑�c���ڷ��ID���!zWlm��į7kO8Q���W��w��t�t1�\cz!�*�Y�i���_[b �r.�K��,}�3u|p4YK�٧:s��$��1Ob/%�Q̤����i�ߺ0�y)褨s.������z��բR��I�	� h�����8�"i�>S�Y�5]H^z��磺��c���&aRTĖcᐢ�T~�0���bW�=S��ҋ��@*t����.d&�ԧ�dwx�k*�9EGtB;�~Y��r@;G2x�!�ݬ
���L�!�!6�C�qT���k�_��dqz �FUPH����P}Z���3�^�+bLvw߯�]o����6�l=�7葁��Dd�>V���/�^����5.�����5�Aߕ{0f#G3�����5��	��F������1��N�B<x���E辶��v �x�e�!�_^^	�ȗx�����x=�CHTe�� )�:z�N�2���D�⼍C���T�^�Bn(���Z/���v/n��2wfo��)R:,J*fǻ��J6$U���g�x�"���	x]� on�̓6��R�ժ���A	�q/�����L��e ���o��c�4�!���VǊfPp�/�t�i���b�$:P�l�`z�y(m����ui_*�x1YM-D���;�,,e�A�f��J���š8�P:jʀ�PKF��.J�i���>��m�7�Γ����gD��Y�ll�tѰ��y���c�J/���?����"	VÓ�p�:�B���<	R4��l����>3/n��@�w�,N,�����@����.�ZQ@ dP����z~��"l�r�/��ԲF��v���)�f p�'?ں��˫Y�Q ����[LMR�}Q��]�ڞt��X�����A=�9��&�A�ZbvV�|Jm\SmS3�}����F;�\���	pإ^s�Fx�?���dp�K��m\��Ia�/����Ǹa�IZzlz�ȡ�� ���vg��� O�#)M����@'�6x���_��b2�����n},��F��
�UCF��k!Hm��,p��L��b:OH8/t�W��g$�&�0��+�.���H�������{?�x�k�B�nx��(|2��8��ݏ�ͷ+���U����%$�^J[)#o��)���$A����/�-��rE����D`(7Ā�|��_bI
��C�Z��hf;`��S�a֤U���R�Ƙa\��jEB9@7PtG�Z���	��T3
��A�% �8KT�5e�d8�0�d/_og=����E��&g��a+�?
�����˜xCdy{w�s4��@�	�e		����E�tvĂ��z=մ��:<��pr�����9�V�{_�#�93��_��b~�[$��蛒�O'����$��cQ�4�B�`�[Ma�����,��u~Ӽ��JZ��qW����t�܁�P|�U�'ٰ�>W�}�T�f�2��]��S=�Y���Ĝ�\�$���🽥,�0x��i�	���-2�3`q�%Y-��W3��W�F��*jq���x��TMe�ӅѶ��&%���-�:��G~\I����PVm)kO�sl��rH�S��Ȟ)�!E]����u&o��p���;R�QO��+�ڪ|�i�1F�bf?�a��V�w�Z�ְ�7�lAn9��T4!\A{��E\8��HS�����h�7@;�\?����A�Sj��XȠj.{
�U6�^�1�N�<�
�`w~R˥�����ؖ�Q҇C�À"�ٻ��3b/��&RF:V�Y��rկ@�c
KB��]�^O&�G��Te�s��@
!-�H������--��~/P�v�U;���'�y�W��y�㊍�m.k
�,����,O0q.帪��P����pS��Б���Ikv���I��y'�G`�6R7��� R.:�iT��u�d�^9ݼd�&.4>�^4�H��8���*e�2^�}�8f*ʷ;���jy4�������<p)���t�mf����SOPX=�?�c�/D��V���7k{YA2
�f�29�_��}Nv�&��~Y�K����M�e����Пөk ng���r5oJN��h:�VG�N֦m[;���O�o���]ɂj"��n�ҞX��0b�d�P�if$�BZLF�R��֯k��v:hr�[�<���aFP��
�������Q\�%�z�{�c��O�)jT��=y��9\� C"��Ӭ�p�c6N��`���E�pJ�2�.[MƤ]��C+���N�z �Z��n��3�>1f�稔<�K���8X�j�o�_�k���DR?vyj���	]eh̆
��^��[i��\�\�n������������N�Q4_�X��J�裳Q�UʈxF薧�L0�y��N��L�C�σ£��3J$٪��y���?�ٽ��"���ڮr�m[o�A� �@y��;]M��Gi.	'9?/�s1�O��O45c��0�
�ͼ�	�`ۛ�Zl6F�ݢ0��I��m׼�q��Ń�,�����(�~�<�O��$P=U�%�)X���?絳��TԾ�Z�2r9�����]oF���f�;���8���߲U+����ҿ�
��������jN�����y���A�y]� w�>��u+�Zgѫ8��6�v�=3/����Ɩ�T"q�����J��=�gZ��{���#^h��x,w�K�ɗ����N�h�[�o��惨�Q)W?r�_1�!Qg�-���O{�,t�.��B'���]�k
�rї�|@�@����W�`&�Z�i����ir�W��1%��tfj�3��}�)	�4��{��v���V�tݖt)V予W���^E�������~�����&���1���U�#�oU��9+t\�dGJ4W�L�2�C=�;Z�6��~�P5ݰw�L7%����s���}4�E��J���է��0Ս��岷kr�/^�ao�A.P=���O{ƽ̦�t��8 K3��!�Q�=�<F0���TR:Ϛ)�E=��td�"q��NG�����n@��rL5�̘�Ç�����`?�]�&uE�a��Ue^�`�M���"7�C�������z� '�l�BBz�M���T�jG�2�	��I���a��]�uq��G7˘	��Jj�ʽ)p��hGh\h��=���Jɀhn	YI>p�2�iK�� $����H\gM+��sZ����ϟD/V�.��ʑBKbb���I���#]kE���>��dY��1ZA��	~�ZJ��7B� l�l}�T����|�tܬ�(��K�W�^�/�"	��$�>g�h�R6؃r�%�0A���u����v� ߵ���g	�<��O�Uu�8q���E8��j�pP��IT/��km� ]�)��4�=K�!�������Ҷ�5����R��?�| _��Y��P����G��؛F�{���&=�P1kl�k�Lݾ�JM.��k3Mw���,b�|e�Y����R�Z`���'�{�l�B���^���C0�Dۧt��t�u��񃣁[���{%��-|+��^������|���-�)i	2���ݽ�=BM1b�:[ս"Ğ�\�U�W��8��;����:fD����q�H�T-�$Ӷ9���Eߟ�"jR�z&�V�|��	��*�'9	��a~�6���'�Yb�ǟ���t,}�v)��([���L��-K��T�Ř!A�9{DU��3��3�K��sɃ���~8�Td��C��>�R��"�����0�︠}s mI��l/h8NIn�E�n�Υx��V�t�#��]���v��=�Bc�f����m�^���=3x$w��bd�.��2��)ZE�9����r.��_S���k4�w�R��`�u�M�wGf��3�I� \Mʾ�b����[�� �r.�|���Ͷ�NAcޘMn6�M�mX�%�f�}!�l�O҉-t�a�:�o���۩��e:NE�n�S.e�}��`u(נ���W�̀��Xg���F+6�\�xnS�&����'���M��A������꺨��;�A���<n�y.ٿp��̀:,o��k�b��ʎmS�)������\;$5�N�RT���.�5CgT+T��P&�q��Ié8�u�j�!$��L��͎�W���'e�~��x�h� I���ׅ�ԎL�-��n�5o1;0�Prʲ�˼I�=�ze_�7�;�L��fa>�P=.i�V�xA������ߓz�8o.�tOw�M����xlP#` \�K�#IR����7�=�7t�`�KA����3�{�(4|Em���M^�$r��ٷ{NPrZ��v%��~�eNc���!1�k�ڐAY�@��-婏�N�����|լP8����x�am�1P���6Q�i�����86�!�64yM���N���F�`�z*3��3�a�H���M���}��G"A�j���㥱��և�y	����d�Ce��Ɂ-@ɸܚ�٭5��`$S��_$��*�a/�l�]9�́l=�}��+O�ي'eD:+���oO�rh\�k~U�w���a�#d��Fr1���6�`'ǆ-���,���*����^�c;f4����a<bҩ^횥>�����]�ǃ���O&�L�ۮ'짴MZ9�w��J�ḿ�+�=�������<)_&��u���A���ʅfj����N�8����3��,���ߙ�*�ه��	���B������ܩb���=�)�$6�:�w\���c*���8��Y�+QW�;�tCE�t����n_�V���������yfe�.L�[F��̏��N��69]�ߖ��3��R�ъ�<n���v�M�F��k-D�a�� ��h0U'�`�c�(�f��4Z)�4�i\��VM}	�Q��aO�L��NúvT�w=ϔb�F�}G��3�PvH	�4���rtg�c�3�]=�Е9BFRgi��IuI�y�8}����L�z��AM���zT0�a�;���!�߶@`w:�Fu�.XX���t;��B�`��w.���5��	n0��Lw%ܕݎ�\)"�/���IRy�n�x��	��T�h����\+{��ţ���ʏb�0u(G�wm�tv��^M��q'	g���'�>XU46�����W��26}j�''[�	v%{��0�m�?M%r����~i`����ܒ69�9�["U朶a��������A+#@�����W��]��O>����:h*4��2v8yumq}y�#,ꁽ����}�$&��L��!��/H
f��@=w�J�p/����l	(��[�y⩳h��9	�q[�M�_����VWZ	��W���?�Fl�����8��6�Ў��V,�p샫D�+����3�7��]�u��QeCzau?�z�#�yA��3�WX=9�!�{,��5�~����.l#��=�c."Q/\�6�T�ã*�����:S2��&�h)��V�wŎsG�n�	��^4Oi��"�����٦}�D�[	{^����63��bp�|<�QcJ�Y�gA]��_.;E<.��y�ȧ�'6JS���RA4$���N�bQ��*Jܡ�U,�\�bwQT���g.8Zl�[��#2�|	�Q�d+I��UXz�kX�����:��t�Q�ś.��t���jIiV��U�ƪk>������q����'$O
�"0��o��v��V��T�p��xl��������(&#P������UP�6{!$|����	g�D���ZV.^r�IӸ�k���e�3����H+�Л���^��7��x^�*f��t�b,?�BP<� �0��;�W�I�*�#}�+�-�ܛh
��k�H�)�5Y���ǃ]�j��>����]�[�L}̮�M3n_K�@�� �Kν��$]�D%�,nR��C��mW��!
�ŋ��ŞGc�}|-G�N��L���R�S��V�kq�mUk��D����Ø���:���l}ھy�2�`��O ��l����٨��?Y��I��cz�*�2�2�L�ǫ��C��2<3�V*�B*KͮX�ɉ�!W .z�g6�z�n��Zd�G����0���ۧ㞪
[zmhb3e��bk�`��U ��:�����W�F/G0�����?@�1ùQ{L�=����#)py�~�>I(��}�fBK����d*Ԉp#�(aǚ��ٚmf���z��{�dLzŴ��f�Hkܟ��P)�Z[��;�6 u&}���F?[�.>{�Z�z"ٶ�n)R�Z�H�<p?��� u�!�h-r@�
I�S�k�8v�Z���x��4Պ���I1ڣԓ`�C5�+l�{�Pb�ʀ��5K���٣irj���wL�O~j�ȓ��&vh6���+�3�e�{r��p3���pe`�s�E��Ҟ���!������^4��I��ܱ���P���oȓ"�@�.na���|9=^d����X����R�.蒆hs���f�1�S�s��!�X��K2{!y���B�G��Si�6&����#s�aF���1w_Ywr
�QC=���e�Z�YDr���o�>j��<%ᮄ�Ǖ���S9��po��FU�k���r���A�8�d�!��-��_�~�^��[�g�lH�c��w`�'�'���)C��/��
�����ZUa6�.A9M�-�D���qܩ�!��؀8_V�x�˒;�2-vwn�����WH�o��] \ݻ�Q����bN����H��Yb)r�)�nF ��D��8g�@(��1��t:~��dR \����OklԘ�>�kAs����;�Ƈ�U�ҕ�����ok@>7!���.�e~&�6��&�:>a�QWԔ��*����첛Ƀ6��Q|��r����2�r����6 ����Ѕ�
%�Y��*6�������'M=-`�y�*>�Ċ{��G�w�L�M'����X�
5K+j��Zlϕ�r�]<��̉�n�F1[�n�6�7Gl?�5��}�W=�4cӂ�ӝ7b��<� ������E����MS3tchvi�$J��$߶�d������خ��瞑�),���^����k�5�e�c$8�N[�P,e�x�/�F�+���@|��	q!���2c�5i���<[�-w�1�*�O���~7k-2[4�|Z���+��x�;�h�6m L���hM����ؼ������2���l�D�#8F����W-Ѳ܈B��+�Gm⓰:�:vI]�	!P2m�d��l`n���Eɹv��=/'7Y����s!^G�!wf	(j���<�1cT�DVs~*��z ,Y��d�6w���ރ�N�G�~h+��C�&�^��7u��o@ބ���\�:�X?�,G�r��z�"�t�
���7�֗Ě�woζV��X��F���vs,�V3����}Nx���ͽ���|�3�� �ֻ�F��'�Q5�7��(whC]Vm�D� l��<�k(�fk����:.PPaQ9p��/xQ�₡/�T���@��W�S���'M���g/w�2Ŷ��<�q5��H�s�����xy�dj{���:{R�إ��ϟX,�^�\��7n&Suɼ�@c��쯿��M6D�B4t4�C�;\^���̈[^w�Qm�5Rl���I�|���ևg��w��Ds�"�2ه.����c?�����6�*�= 72uj�'�)��w74E�w��Z7�<��lڀ��h�=�BL��#{��D²LЩ?�;Y_�I���5���E$�~�"V�ז!�~��W���zǅD�Yih�*�(��P⼻HI�Ȁ6M�w��At1���bh��K]H9��m��@����Ɇ�Av�)#|�~�g��7�y�y��Պ�dA͢�uK��
��GC��9����	�;��u��^�T�X |3��Y�le��A1�D��$���x�w�h~��-R�ԏ�1p��9cW��$�W�Ha�#1�*mN�����9�"�:��g���H�����J96�<0���,����1Di�;T��b1����Pw��S�ʽ�Tt�m�5x�ܲ�K �Զ�dw�S�p%�,��1�d����w���}ص��=��(� o~�Ʒ�X�����S:�P�}�9�¥;j>��Qw��/äSj��G��3?�چv`�Q���̳��g]����d��U�II8H7"�XBL��hG�K�.�
����»�R�{�끛.+�(����u�����%���0����z����X��"���	��s���ޅ���@�֬��Y���z.W*ud�"JH�����;��T��s��EIq��xdpq$��'���gF!a,ⶕ��i��`6�|���r/��T�XB��)�9Fsﱝ�vV�yXDJmW�ɘ��R��,��y,�5�}�qQ/��6���_��ӌՃCu�2^\yC���s_������]ʷi�2(�C� L�3�s��]z���n5Y�ʘ�`m��9�Ō��,�D��>e{XƮ����?:��>X��@�b�,X-$&_׹�M��^�m�Y�+�)�ں�(���֛�P�~��`�M\��
S���q�L�;D����&0ﻍс��2�*,�J'�J�_v�i�ϩ��Θ����w!.yR��P<�����a�a�Q��>^v��h�t��$@����ydt:��l�\6�B�؟f��Ͳ�M�Mm�J��AHA��%](��`T]W�����=��������x�R+���t/_�P*<OׄQ/���Ӣcq��	�k�\s�Q(]��/O�� ��{v��6���QH��5���#J�5�}nns�hN>��f����� �oR�u�,���S<9f�U\A�zH5X��"��]IW��G�q���r6ā@:���M53F+�k�� �q �G��¿	�jSL${'�/a�,�����m�<�.��� ə�ev�жy�A��~�{�1�'�@J��$zf8j�}>�}mlC$�������߲	4��:dg�/78�1F�Zt��S�q]"�jo��g�P��F��(V�%�dmG�C&9��g��	��i7�DV� ���8��y�0b�����@&�	��*"(BljQ�J"A��L��u���
�y�K/������.�Z:�R ������:����Ih�rܭ|���o�po��BJ�,n�q��Nd��tN8��.s�ěj�	��|�[���ݔ"yS�đ�����1/|`�^����5J��)�zȕ��nU��[rt��|g �å�Œ$������YO��v`�t�|�	�}фf˙ѐ�W�_j䛩Q�f�A�P��W�<z+T���E�ӬL^Y�"�X9m@�g�a�n�9�o;�)H]�d����^���ӽ��ts�h~9A��yh��3'��C�:Ѩi,���IVepǰ���8{�Q�������#M�_+a����o� �}�/fhni
�Ѕ�9;Y��M�.��A�?��>}�����R�3y�@M����~����(���t*�w�g6g�q�Ɨ��n���J�.X���x��~����2��4܁^�+D/d`;*�2m��6/|Äڛ����5�7�[�y�g�Ν�T�B����|zK����N�=�b�
����%��I�
��{��[�P~�b.\(���?����A
ږF_��	��^��BS�`Cx.;?g*uʲ˺���$`̨�\p��v�i�u�|�5O~=����C0/���?��a��p��p�Ў�2�=1�4!������w'����l41����4��"��z���W@@�b��GQ�|[ʒ&�/�����U�#O�qPp�c�1�:�:x��w�a�fǩ����J@tmZ~�	�"��t�`�ճ�L!�A!Ш\Cf��U�1�Vs0p=�Jp��ǿ��77�ň`lh��	��(�yKq� *�<�+"$`4�9�Y�%����� $�;���c���G+g��P������{���(���$f<��Xi��U�x�fV�zC�}OO��g�Ewz��s��z���r�dC&)%���	o�*��5�����B�2�@g�-�V�-̍[����)C!���_��v*N��8�Zݶo�<9DH��7!��^j��=�D�ʫ�����3����	#]���s<�[熭#�u*���u����!����3l:��[�`�u�ߖW�*�L���0��T��\N#hX�y�9�4S�j��y�vmi���]$�3�o��z���96�7�lMi0��1<�IP�v�W��Q:Sa$g$z�C /���������b:�����o��E�vqzs�[zq�yqqt
'�)�v=yq�H�	f<?�X���w�e�̤����ߠKɊ��0�l����涩x!���@h=�xEm�n12T?L�l7�@ݫC$��͵Xk�"7V��A�t����ҫ�|��H$�W}�5o/��(4�D��/�]Է'��܂�6`sn�b�:6E�s;��2
+�X�0�������+����bYDt|1-,qA�w��G=����T\UO�h$��=�x�=NԄ5:�i���$�n�A+G��r<.�׏6�8�	7Q���� V n�����%��C�r�7s������:���>Y�w{s�G{"��?fD�֢	��c5��Ɏ̴�yҐm�Ğ�(\�ȁz\��[w�W~��s߮DpB�Ƴ"����</U\��yJ%΀�4ϱY$ᕫ,�U��;�����<�Ϗ���A� ���(��@�ܻ� �{e?"�fxc�[ &s�d=��2������!u�\c��n�D��b�&j_󒎢J&�)�T���h"yN�j�j�y
p~XU�j��J�p�=�������∻�Čx��Ⱥ�}x���s5x�2�V#�d�ضt�� e?ͭ���{���33j��-f����go��Ab��$�-��:��lAP/=_٫����5&<��!�T�Ēg��ċi,U>E�<?���lV��#�����q���L�]�t�����	����GLbQ�#$�|mx��w�r\�]"�B��(jrCY��N�SUG�ٴ[���E�9��C���-m��*d����������5��+EL�ȭD7>x�-�6[��'B
���Q���~�[��F��;'��0���G~[ꖺ��F��rc����J�<J�n�7t����/��h��p��~�l���$��[�+&;P�\�p�{ɩB�p&χ�Iv�b��)�����D/�h�B#+�z�!z-6ej�Ɨ�a���+�|��M]ϕ�Td���m���{>**a��Yt¦ƻ�GNl1m�������}afT`��b4"��ިt_Z��E��F�hP�����o�$#�E��p;G�<�"�ˀ,(T�|7M]���B�d<�!TBw >_K�w6�����G�}:�_�Q��陛�:pM�5��֡�t�WӸ]9zc+����b�&q��=�a����"�cJ�l�|D��
vWzI���w� oО½J����e¬� g�y}3gJ�Q�3z�eu@�'�ufS��K<�e2n(�ojT��d���Ѹ�����ر�
5��b��6'k�V�@�׼)`�4MJ�9�y�0��>}��n�/ҕ�ɰ�\̠��/	W�fy��W��7\s:�����cP(���R%`g{e!T���w,<���I�2il��[ 4�y~m�>pF�U�����s��V_�GI���?!��o�A��JD�-��mk4T��<����k(e��0��	�g�d`-��L�" ��yg2/SQ1d�<�(����}�L���;Zb����{i��Y:��[wy/������#��|�����F�q�$��qu;����gDV�:/ܽ�"�N�a	?p�B�%ֺq�R-��r2	��	�V1!���S���� /�[B%�"�uM7��f���r`r���x�BՏ��[�wjtv��J���&a�����{sL�3I��Z���m�1"��-���p�(O�b�@��/J<��0��}�^�j�׍�82%qs����DIh��v����(���T�x�N
Y(X��b���V��l�7W��8SK����!{wAh^���!��ʾ.H@��ٖ����2�XxX�P��o��1��^�՝^:�������.A�`�
r43�bJ�i�=8�<��g� ��
:j��y,(���=9:5�X(e�^F�4䩏y�u�[A�.�Ra�W�Q�̐"�v�o���s��K�Yk�����ENZ5���i~x��Q�z8xޛu�^FLǰ�6���yQ ck;P�J�]Ƭ/%�KE;�.6��Q߼޾�	`U��Ǡd��ujy_#�O����ٜ����eg�O5��0��������MCT�JM��b��e-X�.X2�w�C���v3"g������P��f�n�NsQ
(����z��n�q�/MG��o��j�!$�ŵ�_K^���7���! 0+�Rd�%Hc$i� ��~�ӂ�x�˥�B�v�}�ճB��ߴ��̗q��V�Y��F�V�o�p�[�g#��^�;�XhC��hv��D?� WSwj�b���I$���G��`������Q��C]"{���	�>_��W�5!9b�{�a���z(�
%.E�snNԨ�p8�����G>��b`��e� =#��oY�O�tҡ��﹛�]�斡b�V�>:v��\���ے�VI�=�M���d{'f�6�� r�]_3q� �d+XAB��A�pm�G�L�?ʝϓC�|����;�>I��d�^���`��|�+����xu-/�f�"�''�	��/<a;��ӤU
�!s.�y�~�V3t�&N�δ�����kL����K��{�:����o��h�ci�ڡj������5W�ԠQ�W�r��|�nXK�wh��tֈ9��O�@��L��D�zI��᠍�>� z��8�i��jpƨ-.�'�5�r�r��k�M�ґ~v���H�1�Z8�S� �ON z �;�Ӳ�o+}C��|�-���!guK/&�I���.��x��s���2n&U?yO5�E�)���1���Y�mշ�U.�����g��M`{_R�Yڥwp%�Of�5�v1i�vst��!U�|5�:M�� T��ɦҀd��E���z,���� �"���<�We_yB�o=Eٌ���ߝ���2W4��_���E4�b����4�z�Yl.dJ��9&��i�P�Z�G��4�>�lYMЭ���/�a����Y�K �[f�룬���XB-���/��{�2�`[7�&��u՘��st�����F��?�S��0���lF�st�����䯔��U ��EƊ\�$V�����{vO���r�省$�u�Up�d�%+��3 �����Y�`5��Z5��O3
�B	�ϝ��H8�B����1m'e�$�����Z�ooL'Hu�jx�PL^L%�cgT��D<�Z)�;ϕ����M.c����b3qPD�#�nξ<1e�b�\��=�hA?ĳ��t~ �����H�^&�����0�GX�Mc�*n>���'�m�{C�ew�:���\��2�,Rݝ��1�����`�4M���(t>S�}�*�]r>��0i���XH>������Y�H���2ŕ��ߵM��v�Cd$CC.��q���[P(����vj�
a����ա돆*y�Q�|���YOv�&�IY J"'�ձ}&���wd�~�k��� �r����UN�c2ДL+��Ɉ6M�P�� �$����g��(�9U5�?���}�����E�ӻ2l�;�\Z�ѡ�_�m��[Թ���-7��ٲt�jm��d��D����rҐ�V�=x���VA[�}�ᄞ!�{(r�ыn������{�p4��A���<$��ߗ���i��A��l�Q�Y�tx�U���A���O~�]i�yu�i[���/A��ސ��+x�G:���뫆�Ȣ����N G�w�]�Y�͍<�KT�������B��e�\���nx~V�
zE�N�-�*5O.�% x)x�WϘ��XdC����؀ꔳ3 �Q7�|����ۡ���n�q~Hje�A�R��}^�]� 8�7��=k��s�����X��Sч:[]i�9:�i��9Zr9��tʸ���.��c����&���|�'_��n�����]`�L Xe�,N	O�I�c�=0�M&�Q�h_/����a�-�v8.�e���Mݟ4����ߛvlC�;���)�7��|�� T�Z��D�u����F��MOԖV��t}oe���+ [���/C5��Â�Ż!�(�yEp5v�^��	���dB�Wm3)��[�`���r�
S��3�
o���G�-`|W�j?��i2.��p
M�u�f4z�F��9s:��(Λ�Y^o�E+��7�kX�w'��'�� $-P�
Ě@e����%�;���a��,¢�1`��#��Cy�O��4��H�#i1h9�*lJ�?*�=�)N1=�1%�� �2���hc��d�����3Nti�ź8��&���a7�{RZ(�Y���B���$N��PY�/X/�g�����vO���� ��ƎHXoq�~bL���(�-K�������.E�pQ�'J���p)!�>��KҍY��.ݢ��Y$����'$z��������=��KU�n��~	�_��y���Jt�K��v;��!�/#��;��TF<��q�|��`���X�>�	K٧�k�Ed������j�c� Ջ�]����∷΀�t.��"C�a�M�*�;�6*-1@���������H��(�����]�^k&��(]��������H�$J���uD�
ւf����M=�7(��̶��nb|�y�Ʈ��-=�$jb1eq�؈ǝ�)��O�|ya�2�p��n�3���Q^N������ň=n�=\�
���
�R�J?�x�G}m����T�tAaG\|�����[,�U;��Q��{s�?�<C�I���}�&���D@E�b?�����`/}3�8�EiiT��H�&	4SO:��=_�[������>�6��1?]7B�i��yC�h�O~���UZ��ʹ��q5��:�p��U������YQ=���s`� umg~[:_��d4evOnI�Y���ro��(�$��{����U�ǵ.�B���<�g��[y��`ӵ֒�Z(+(�@tN\�:�1�ŀk�*�nuy���6.�k$�?�Z�c�sKZ��pR�������Ns#;�h=r��mC���y��/�X����(.��^Tv�.p�g�b��⚛�"���L޳C���Ps��
4w;(��jvB^�`�K�gkΟ�yi뗒�S/m:�7j0��X7�����z偾a�nq������tW�Z�  ߐ��4�@r� m_���^R�~�s�@�8��̓�up�A.�Z�;����o�ֱ������^�m�
�c�����]�)�/"��/��6�>����}D�d��T�v���C���,i�KG=W��ٌ=-o1c�\� 9�3��O�G{� ���;A�J$����ڲV�s�q�	�]F��v&�Կ��-돋�F?{}yZl��!�o���[X�1�V�"��_P�F��/fZ>-�pPÞ_ J9SE& �k��
"z��P޸��2������H18b<�cx��w���m}%�G����{��K˯ҝ�l��S�b��HZ"��O	=�2��-����� �I^�C�7�Dx8~��:���*��~YI�:�ݘ��:*��}�o�#�J*W�"䰬�S�։J�+r�v��Y���:����b��VElΟXE>
�93@ !��m.s�GtS��(�P��G]<�UBI] K�����z]���#��o�ZٌN����]�e�����8�����s���m�V6\�$ţDU̶�k!l�&����9O�����W�Yb~x�?�{���	r�7/�(����A�OJ���2���B�j�>(Pp�3���OR��>�sn�Wr���CA�@0���$�OFn�@r���0�u��"I�Ä3�]��w�\h�����²	:��#�?*tVw�sg����gj��o����>��ϊ��q���lgMp��ȇ��(�dn�w�Z�k��
?ע�T4lyT����0`��x>I�t��N��Jwe�t^!��L<(�sۏt:�&+ؼ��� �3�Π�%d���4�@���Lu�NQ���V�s.��Nu��Y�v�s��
�������c2�f�{y�i
G��:S�B�B�,����n��G�g��&��Iůd.�/?�Ldk�h�y^�1��$�<�a�ִ�=�Y��2�~��p跜� !+/��Y�ud4E�n�2���/s�+.��ȕ)�S~���S=�f+�$��E�ꝴ���k�����DI	�p�*�,%��ּ����ͩA`�Hz�FE!|d�̰�J#B�L�OWy4e bL�Zn�Ι�|L+�Xm����U-�'{U�+%���Ӱ&��Y����������$"'�X�@$O9f���W�}%.����:lz:K�v�F.by?V��ؗ�],�@y���nK��I�p<L��qv��B�l��ܘx��QKȴj�y���� #9�-�+�S��?��[��w1뗅�q����8W�	%�u���ْā\�
�N��.���Cܨ��o� �Q����Z�����pua��	�5پ�a(�K"�W�F�y#�;|NnZ�$>2GC=� ��8���6K��Bi�ь�x�x`9��«�������)�_'e,����b�6���7�4�z����E���<��_{ ��h��
i���Q�l;o�%�uEQ1�v��A�����h����[+��6	P��CC�'!�����j��85�U��\C���B:�AOR��}�f$\As3FM����V�� O��X�塙tc�S=�%�Kت������넛��㑕	a�Ҹ��oKi.E�K�m�_�<��G!�B�/���OQ��4���9��.+ѣ��Av��:@8��
��n�f��)�X���j�$�)��j�c�ll5�8�7��b=ֵ�ؕe�brOo�-B����(B�9��q?�
�T,�W��0�VK�3���]Ij���V����"�������*�H�<4y���V)g׵qz�0�ѳ��'�s^�H�񨻜.������,������~�����o� ���r���<�+��|��������|�ᇗ��?߅!�~������zJү�����T�3E�N��Z�A��Z�E��e��3z��Vi��q�E����p�WgfAn��z���.������)�$��p�����ͯo-��"PU&{dp'�O�*��U'^��%;�^�]����\86j�]�@����"X�J{�������s-:��1�0�	�`�h�#��ݒFq�"3N����	ʽ��V�^�:xS�o5��N�v�A�,f�t���6��j��ٹ����rL���%u��С	�ȇW�x�t�' ��7�1m	�ikl=�i�2�2"䷄ZK_C7A������%��E��PqA����p��(i4�X��1u_m}Pw+Y��~���
����������9J'%���������C�{��͝�M�_���M�,�Eq}�怖8���,\����S:%���
���r�*���"�ě1n���9�G����;$E35��.�.��H�e���|���p�h�ϴVP&[��G�H�"<�݈�s��I�G��ແ+H<J�@ky1?+D�?2Gd�9���|^�[�U����G}ayR�#mT�Ry��ѩzS�3��䔼A�&gK�z^[�2u��w� �g���&Źs��Y�`�=>���P�wDА���D�5Q-l{�U�\d��@-�\��9��� -T�K;c��yVԘ;k�Q�?/v<�Ƀz�h����%C�C�'ܘ�(g���Ĺ�-�FmW�{�<�tnM��ߎ[��f���^���$F�5N=\�Gn\_>���b�/���N��%���	%p�]K��w�A����r�p�%C�y^N]ĢB� �q��]�k_�{��,e[�Q���ƙ���ˊP�m����#u:ok1XW���B:ԭ��M��0,�����6�� 1Vq��䩉�zU(���� u� �gl='���7��M4�O�(�O���p�Q�v+����$��C;�'�w0;C`]Ƀ���7�)BV���6��0B|��2C���3�K%�\j������1��8Z#�G_z���=1�S�����(S�w�C��.v��_ʸ�ޓ�T4�bN�]�_� ���8u%<]�S ɢCI��K�9Yx��N-/�6фK(u����PmS"o��s���ŐV1t�\8��~ɼJ�P>�z��ݤ���g��[�(U����eG�k<e���ӆK�E�� ͖�ƥkufm���ҔK���tQ�����zW��E���6G�N>bXYc���4R��o�%i�����	����s�J��!��X�0���v�!����Ur�Ѝ׵�XD�R��� 9nM7����ں�4�k� 0���C�n9p8��L�j�Z������g��v�3]�gI�x_�X�qgΔ$���i������'�W	X'r��էBcZ�_-���7���쨡���kv����#4F�!��w��D��������9��Ԇݭ{R�?lU���Q4\��O�݈��Q'QO����RE�/�sa���d���?���OAJ�@��Uv��%�v���V�a@ ���fP�w�������Й��ʲ��uL�_�t��-4QI�X�w$����õf⠶�������խ��̞*�MY[�3�l �sO��]'���qҥ�}o	��\��Ҁ�f�C�/�x��A�X�p�B5Y���FƕL�>q7��%-��}5h3�|��,���1#i��1�h#�@/�6\��ޕ��d�V�[�ȧ�!���8i���]
A�B��QC������֐*�O�u��"4���(��VQ�sR}Ƚ����u����/�8�L�t��cs�
�o�f��:eGg�L^�N���Y�#.yH/�G�@b��'�y��b@��b!�1��("������A����2!
9���bL�N�.����q�s�I[�G;SN� ����2�g�XG_�O~p�l�ZoKqA#`]Y���|�t�#�iZ��X��:b�B>D8.�Q^���^��o�����4��qW�gÇ�P�F�����hLt
wV���{��n<w�J���o�����0������� +�>�FK��j�ZO�h0�t�����PΟU5:/1	q3N��Av{�?�l�26��,�k]�Ę�������||W����N }��D���5
�!F
��hB�h��بy�cU=nA�S?���;�t:o�e�pId�E��0���'���֬�r��s	̋w��h��Y��4R�mN(8�7>���*�
��K��*����-JA��&p����Rx�t�%<yr�6�z=#�7�b�����0��.��A7[���ۀ�/@����j8l�Yj1� \���-����x��6�C*;�Ҙ������'��Rh�<�
n=J��U��f�49�ÚE���#!����æ���h�=���F2垦̙�s6���ǉ$c�gYFY:��P.���������RS#� V��d_��D�]� AQ�-q@�
���U_5���T��H5$a
�!W�&��q��m�Z�M��TT��Ǘ�G"b�����D4�5��=^�8r��
��B/��T�ZuWd��#@��
yP���o�n�H�1D�� �]��Nb�F�2U!Pu��Ì�%�g�z�:�#9�!�[��7��O��u�r��{J��o�QcW� �Pp{�D>�0,��'▒���h�
�Qr�y��Q�G)i�%��W���+ޚ�s��^�L����ɯ�~3b�NCA�e��y�=؍�a� ���d+�����"��?�}*?�ٕ5SBQ�r4rR^�y�e�:��?�8 �ӄǨQ'6�g�,.���.�@��J^�魺���)�uղ�����K/jð0�f��2���(��@�x�ؾp���aO�	3Es��M�Aj1?	�"�*�y¯y��1�$H�g$K^O���ӆ���r��,�?iI#iDZq+Π���"���=�}�( �q��7[���i���[�)#G ���Ze�����#M���x&?Q!K���ty+��3��)C�՛̼�����*#E�cg1��p�m/,���Sw��hT9=Jk��/5w���|�@N��Y�#	6���J���;�e��Go���
��"�k�<�q�C�.�9��6jS��U&;%*uv��ON!�jV��paO"�Q��$}q���ط��3��㎂�	v���ƛ鲙٤��\Cf�c��7^{,=�RY4�8���hu�^�`�PUŰ�-���*t.�Y��A�����AO��Sb���ԴBr�.TH�X������I`��
V"ϣ�8r�;�/��p�fKq(FPq���	dY�?˫9,�GD/�6�ɡ��Z��{�$�p&l&��6����%�.&엧�1xB���v��"���s�X{�˅�B�@�
<�O�,(��F7�����f�7J�me�6'=�>��,X���r�r?�H�r���coO�$���+�gH׎�~�1�|Q-J�Ny�g��
E��r���#�����gBn���+���=q;��6�S^�6��>��ҵP7
�0�0>s���<�����䫀���p@��ol	��O,��sr%�D�dJ�Z���r�ʠ8Ç������>�ϼ	��O���`M&�(�T���rvCPn@Vo�</l���h���ti��!�3A{�A��x� R9K�A�dnNK	�ç�9*Mk���E>��>V�"i���VCz�i;7}AF{��iAƸ[�ʃ$���<+֒%G\��1Q8�]z���_3# �P��S����d�d��)�&�Aj���	��ҍ%�v�B}d@���Q��a�b;��#��2,E��̰{����U���ay�}�-�I@�#����|<>�K��5����h&����Dfv�	������r�. �xJ�hC���a�ԗ��إ�O�h�CGGA�n�1
�.�ud^��1����!O��sB�K��L����g["~���"�����V�g�D>�臘'�ob<����e)��{9.��m
��+�tm�̝�rRbE%���S���&]�7��Yb;pGs���K&z��\�U�����r ~�.�,�-t�@�-���4�{�Ab)A���mR,�`Է�	���.sm��=�T��n�����Ѕ9�+#��b��[ۍ6����&ʿtL��&�� ~�<�94��Χ���=�fʏ6=D�2-|�|x�����X�m8����]a�Z8�2F��M�>Ӵ��AL��^K�zEv$/��)���f����߆!�49(6"����R=�f���+&�2��1�]�.b*k{�}��S�}�Fo������ �,���`�	��n�J[�ʣN����mz�������}�Q8o��������qߵc�h}�"N�xX �B���[�~mSM�p#�l����_D)����jd+'��o:�9ZG��C��N��m��O�j��)����@�BQ��[-ݧP��λÐP�I�X$�u�t���u�q��ҽ�d��<�^n�d5P��31���45ǅ�@��rvHb
�[�5�D( 	|u@:���֧�dg}s���@'U,����'����FF�0����0���}����M��OW���Sʷ����5���c�U�W;�(������.���z�)�,n�[���DKm��5��~��3^cf)J!������"�Z���Ǩ%$Ȥ���G5�|G%d�!պ�ڜz���/ T�PgL˷�{MI]b�<�G��G��@���w>QIY��u/���B�S_wJ
�׹O`��"��<��GQ���(�ED:�����@�����I�<��H/���TX�^��F������|�\��z�BɞVIb���V��ŀ�K��jnΞ�CZpF	hx�1K`Bߟ�"]�8���Dq�$�\4?�����a�GV�O�(���"�H�ƶ�h���o�9s�c��E�T'|�*p�y�bb"�>f�F{\�1�sɐp ��#���I)Yd"(L����C�#�e(m�j�0p����Eu�J4�Aun�?�׵��w6O^S�)t�^�<�+�� ��hŋ>zЙ��Z˰�iM"R�'�� �?�4�}a�M�����3���@���B�-��7�N��b��m��fv_q��ȗ	Z����9���	M�e�UJ��^��̍�v��iV��4���h7b��V���U�4���GK^��8����� \V�fS�׃��D�a�x����#[���X��q)}���ζ[�8
�p�X��pe(��+�{����O�j	�ǯL�tJS`�P�x��(�9M��avMcv�ytp�ܾ�/�U��NVP>�wbw��ZC�
�=/�ע�=�h�9�eve����[���6vJ��1���)?,��s��UΤ�Eߧ�i2�uxq�6��,�ܨo��>��f�3��>1�؏ٸ�[�o�DJ� ���`Tm��S�v�|�X��?�)� �:���g��xd�j6��?i&ߨ3?}�ˆ���-"�kP��_<Cs��-�֛]:���6b/��ڊ�n��ح�_���ɇ �tCN���X�WOX��{9
��D~y$Wh��#P�c�&w�8���,�R$O��!����J���}c_� (|�R�V�MZ�o�:Pt� }5&݄�q��k8�� �c�� �8u.�hFUU:[�����t�}S1yp{�d�@���ĭ\ڗK����4�Q����l�φ����,v��M���{���G.���`8��Ys�2��Y�ֻ'�5����c��^	O��k�"�c�#wx���R ^Xɓ0�����);0	H$���$?/A����ҫ_������-N��IbG�|�h�4�i���ߞzr�.��~�y�E����>q��.��L����ٷy��!DS��_����lUf7���5?&��ȕ�	�r�Ϩ5n��ݡ��'��_n�Xx�k�g)��-9�zr�]f�-M���+Hiq#+��&@ Q�\��͊n5���?�q��l��ݳ��S��8!�q],�ip�o��oQ`Ol����m��R�H{4�Y*�|��`��E9��*���|�IcO`��B��s�(��N]N �� ���T���)���82��z?�MA$�[Ȑ�hS����t��s�@��$=n��p�P�kq�!$�ii�$i�L�ht.�1^�hVRρ��pK�GA@P� ��#{�o?:^3V>�/���@�"�����D�GCo�w�6e��"����2������������u�"d{F�s5xN���X亾� #W��� �`�����<I�w�տYK�
F��Y�H6qO�h�UŴJ� �qߐ��6��/�X�z{5����I\��x>rc?��
0	C�����ˢ�
��_��ٖ��b�b�m�v���F��3��������4�.!�1O���G��w����޼�ˉ�K�&�)v���s�-�z�束������nN>��W��5��t��Tf���1�n��؎_�E�P�+�c'K�<�m.�2*&2��EC�j­��c_��*�&��_�"�>��Z4��4��9���Py�CA�?��E��@�l/�6s�W��\0ķ.bW:_����t�n�ǖ�=�1t�����F��c
��RzE������!�)�P�L!���L�)*�5 �fbc> $�||����7�ê֜z�n:ӂє��i��/�~�J*�m-jϼ#������϶<��dggi6	�4�w�Y���`$���%��9�ZWz�-ˁ> ��?�p+-՗����lZJ�8M�8��m4�d��v`4�d�<�\a�ٞ�>.蹈�f��Î�8��hu��m��z&Hem�		)�A%Ǡ���GR���=��S�Wm��14P�/���^����jݧ�O��j����� Q�ZSSߨ����9B:��l����P��`�*���:��k|��[�ѐ�HwXL�[���7�f�D�>U.�JdS��HVu�}�Ej;�BO�����i�����X�TQ�L��ľt�E%m��AL�f:�o�{���0�V�h΋w�"�!P�?V���<�E}�F�]'q���#x�����OZse�/d��͏���>��
�
�R�	9���6�&�g+8�8�f�H�UTrN B����_IF~�uAשE�����e�'�5���X8Bh�(
���&ڞ����̄��#��&�x��5�,����z�S9���EJ�a'�{���g�{GG��y%�:�����o&�[_K3�SgRG#�vԿZR�������3���7��6+�#Ҹ���� ��wvԕ��Q�����Mm�ZwaIZ��H]ă�EB̢�G�`��uJ����;v��|�t���m�)`�!���9\�<hH)s8�;�� 6#�?=rs����ʑJ��Knݏ�F�u<(���!1�h������|)x�:ro:o/T}���%`9"t��&$1�����h$}4�Cڍ5w`a��l�2J1����[�Z�����aM�������5QȽ�0�}�FZi��?jY�(��8�O��L�Q�#@쨭������!0W��sCXh�3Z%�l�I�xs������J�u#�EU���]*4���%��$���R���j�~��,ix�k[헙NF��`�� S�U��뀞�4��7+�
�1���$W����B��~%n���vdp~��dL&�Ȱ�M�,�(K'�� ���V���m4�6�yw��6��̀����.�C�]�e��DEЊC�EǷ+�-��\�h��(}Q�9���t����)ne�B���W�Ze_�A˿��� ��F���0
=��T�X��q��ץI��}�i�by�����Ez��N�I/ߋ\�ʾhc�L��7�~htA�3��p�����>���)��_��;�?��+K@�N��ǵ�w�
�0�*����'�$�׊�*-��޾x]�n�D�k���S^:��"b��Pes�̖6�f�&�L�-@�
�0N��!��/���kIb9�7'g�H����8��B�r9_�+j�w7
1���a�}2mcÃ��S��xL�E�A� K4P ���ߐ��sTd~�aa��y��2��M��Id����r?ȥ�!� ����u���`F͖�IQ�9F��V�P%9�w�3>\f������̥��g���#���1�ỉļ���r%L�#}gn�@2�W�c��?�D"h$���F�SW��&g��꡹�dn[I���BF@S�K]��m�E��I��;%�ᔧ�xqݰ����'?����y�|g�n|��C`���	���c�s0�3$x7?�1�}c��^�#J�ƶe�xtN�x�kP<�Jl@+<��Je�t-�n�iq�~w��Bt��u��m^�u�O{�"vXU,�e.z�+�6P#�.b� ��\�&ρ����v��#�!� 7�8_�>oW�jsB����w9bM�X��P��ǠmkxQ���r6�km�hH�P��þʍ�)�g�W��=�;~�F��i���eծ�o�:�����6]�h�cs��n��DfTb�H�Zxw�LYat�j~��g5�ءvt�t���h4D��Q��C�ne<�=6�K�9xd�Ꝁ�pfp�7�Z�&��LlK�������A��3�o�\��}%�ɒ_��[_�0c�k��^85��:�5@$Z�6^�D�N������p:���B��{��}��BZZ}�NvpL��wn���,��e:��ƀH����I�>5!O'��H��L��jO�}"{�|ɉ��Ob��	|j�� �z������b��B`�.h�Y+���\�LE��K�S�[�����q��E��Dܜ1]z�����cأ��a~���g)h�P��AA+h���d��įĤwi.
E�"�_����R�L��P�xz�R}��?p���l��8��m튙������k�z-D(�	�4k#�(�b��
�X#)�!5;�Q�&��iNT/��0G��L��i�XΗӸ�z9�eF����2+:�w�q�>��|�Q?��!l.U���@7����[���q�w��t|�������ڬM�К��طg�Qz[��g���A3�����=]�
l~�'�k��1h�q]�U���'��bM����Ѣ�!���^�e��2�r�ȹ�;�Za�c86�`(V�^=����ʌ,�XJF�xj��3��IZϩ��3�mm�cԛj�!)���8�O���V��'��!E��֊.E�z�j�BV&T�1�.��Z"xv��[9w��YL������D��]HMD�&^�I>x�s�u���inN��Tƴ�tp��|�5i����촪lM�<ᨾ��m1�t���������_��G��=�eZ���U�+ZIu��	�O���׭|h�@[�
���v�d)e]U�_���q��.8�;9���	 �Ϙ�8�N��1ӎ�谸3�)
�81.�.[��9�P]��yn�J��[q�lP�%b����\v�lK�7
��/K�����CO���^�g�S�]Ӳ�{J�(�:�;p8C��6��p���f6�G����������J�1�w���<w	� �MP�9&�
g}�N�3�ZZ���C�8i
���'�ٚZc�Up!��44GY�������,��vK�;;����h�"&%�NaG�v�/:2	��(Q��E~~�c�]�¬��!��-�J�n6�?v��go��gXG)c�O��F�j {ʠ�Ϊs��kШ+�:�0������9<ў$3�sZ/3ע�g��^ʙ�2��mU��Z��]��%��-��v1������qC��A8���@ǐ�D�6����Ȥ#��*�L�N�E�;|�m87���u��Nk���D<���_/|
;���Ūz��a��m�F���3k�l����iv�����y�:���N(�w�k�Q�ȓ<ؕ��]�0m%b���#���S)��JL*�w��,?��̰R��1{s���CB��<,�� l����Կ:=e��9:�����QF��%X~=;��U1m�k�7���T�/eWg-/��}�"Y�q�Z�<I[��]�WU���vڧb���U�IH��Tv�,���fhs��N���+�r��'ݯ���5Y~<�ma��jW b�7�d���-�ڢ��\3}\\ k,��G����E��#xl|�{�r4��G�ia훉46�?MN�ܔ]��)h&c��z�XU����X� ���g����ۭ��r��
t��!5�x���7|I-'��2p�S6�cB����
>k�o��򄰥�w����c#q�;+�(ӛ�k߆�^	������� E����~�Q�e=��J1%�Sy�5����������s7����AY5�u-x�8� zW!|�C"�<\qHU���|�	K-���ƋudM�T���|Jk��k�1'�M�F#�ĵ?";�8&�-�,��豢*�N�ɚR���M���b��m]s��a����'G��P?�ht��dڻ�P����
fw�R;�t�V_;�3
�S�bFxGZ���cSӢ�>j"%
*R�3��v[e4jBUΉ�
�j�!C9���������9�hM�T���rDfJ\���[�u@K��7&�4�htc��a���ɍ7�qhԘ�/.���O�_�,l��{���% UA$��ay��Ʈ=�Se@<W0ϊ(I	����y���!+m��y�!Cc��A=d���:Z�Ue�~V��j�:�m�#�0�,i$�D�����?H\�R<�����9�[�YG/fA�O+����G�_���BF�@�&0��X�ϐ�t�[P����f/��`u>��
���c(֫�6:I�v�����:��@��D(�(��~�8�Ѽ(�Q�ӛxƆ�{��뙤��2B�9����3^n.�=����֌���d��_Q[up��i��{3z)� ��ؒ콖`��r�w�.c��f�>B�*\��p�_�Ɉ2�|�f�i����Κ�ė�z�8`��ƣ������>+uhn��m��5Ov�+T�q.̐φJ����/����C�4���Ҋ�t���usw�,�ΊX6CC���������
�X\���#��s��'��u�4n�RI
������Ln�Uyr߄c�x�?oIӑJ����_I�!^F�JƁ��\�X��rܴ�TmS�K���ʔ?��8Y=��f�t�Sb��fJ$��G�֬��_�\�y���_�ٺ^��&�n�Ըuhϴ�@��4U_נ+��|8����lb"��i�?1e962	oю�m��b�/e����1�g��%��!L"��di�����âDf��O�E@+�2���o	��ys�&n�d���W��i��}M��W1�.�s���J����,kI���G�����o���vΠ"���n;���e#�ȽZ�҂��)t���B�ׂJp|k��~���qU&Z�����ɟ����iO��	��c���CWf��Xۛ��$]�_y��d��g �q�c�uMh�rb���]	&��h\��?������y���e~b��x<uA2�IVO	�$x�Ǽ��������L�s|��Y�bNa��H�0�F���Ή�r��#du�s�'/�g^<�K&����cJ;��4olUK��k�ϼ�'�
cD���#MAV&Q�@��~�1 � xM9`�>��y���t����/��bk�Œek͠��k�a�A�n����r`+���څ˓��>I�߁��	���r�wt�
m|�,��� U|
8�Yʖ��5��gUp�@�)���Jg�����+5�Z
uՠe�8O�n�4�)��f��-׀@��m����g�����I'����-�$#���I.�V�`�1[a�4	���Q��m������{%���$L���7�m�z� ����^]�;�z�ۻj���Y���֝�O�dx��Ц��:!�2�+Yi�wY}�����:�Pa{���'n�:T@����96�j�'yN`Q�4��y�Tw+L�j�1�+�`�<�Q�B���7ξ(@�Z��g�<�jO"B8=mPʭd��Z/�J���B}7q1�,Y�Q��l�v��Q@8�C�7�yZ� ~~���y�������*��=}������0���_����\���dф�=ULn}$i�stY�|�`s�̖,\��AMHt{G�(��{~˸��e2�j���V)���T#4ڱ��`�[\�6z���hR��y�/%��uD��`!�����(�om7�	&�|�0<�{;C��[]d��z��b��k�(��%��2������hJ�w�?�����[�ߥ�z*ZG9B�	�=�[������(�%����:���kAW��;�ZSՉ5_ܽ$֭G\��X��51,]>H����0`��P��������(,(X~[U�X�@�s��[���w�l�
��/�9O	,>z����V���)�lw.4	�kY��IA��킋۟��������	�^��q����.����Ӂ,�q�c�Jl��I(yt/�F@�}~��jZ� Y6�J�$�bGa&�iH��'�a�S�]���(ϊ4>�I��$m��i�[������k�JM}�m��k��W�����3�'�w�u��D���bB%��^#����Џe}��!��j�	���A��*.1�2+臧�RZ1�u�X"squ	�
G�PԠۑߚw�z�I�ƛ�D�+���j�v���A��G�J��Q�Y�	��N�G*Pa��wZ� U���/̆R!�x����Lɻ�	2y��"��S��^u\BZ	��tKUi(�Ζ-$�3)��ۜx�%���=�l`����`ȇ�}̷�K6]T���Y3+�h��3��E�-�gğ¼{�٣Ϙʲ[e�Z�\�Yw��msiϣ���[W�aİM�{�FD��0�,t�Wx�4X����p��=��0G�G�>l�0�0�yH�����,�E'ϰ�
P�=��\����Q��x���[��_�l�3G���Z����_��f�+D^) /����J�Y/�-n���W�ÍE�U����~&��?�a�� 1)�t�Q�2h�{L����v�̞� ��A�M��*讂_��ȮV�GG�;	���7��I���%����@�{�TM~��^�%�J�
�a���uz�X��6Aq���z7)^n�e��3I��|���1ZJ�L=p�&��� �'i���j%Qs������M!d��\d��j���G�u�D�G���&����h��Gf��.����Y���pw��ݘ�D��><�8Gsw�Z��7�*$�f�F��R��"��DKXoy[��+�m����*Nx��CR+�,��]����[������t[D�m���lW�������$�iPW}��B_�`@Hd_~�\W��v*K �쀚N|�` �x	��P\��b%��Y+B������c�K�����BZ�b���L7�$I���������AOv�ͽ2��H,>�U�J����V���J��$Il����%m�ɧ���/ԗC��=���+�"�
��Q�~B]
�r��p�O���(��a58%8d;�-,������e��_Е�X("Md���s5n��j�0�G>�;C��αj��ڮ$g��w��UR�!�[��8b�=�&Ē������0�iHS�L�g�)!b�]Km���}�z96C�Ɵ�]G���b�0�N�K?�3�;�b�4��-PH�[�=/C�M�'�����_x�bRjzvz�&L�r�t�{�P�m������4�e��p3*��EV�n�de|����;ļ8n'�ϲ����E�$�q&:9�툾���I��>q�Ux�u3䕑��Y;��9g�����n �k�������i@�=m��,ܬ�W��^��``�,��ʮK�a0�.ݎ�<�N�#?s6&�)be��$ �&�d���=\v^��jDI{� ����2�� ��!����$,E��ZZ���o�W�; p�F�@�s��-�?��&���;o����������I��\B�Ng�8^/��a\
��6S��$���2��8c�R���6��yB�'�
�L�\3�tג+���I!2�|��|ZFW���@�����~��A�,�	�[��=̉�\;��$�"�:-�D^`�ݙV�T(��;�џ�����Ay-����S5�0|�Pc��m��W��!�Z�wЪ�)I23���K����!��Y|��BR���x��T���ꏵKʁ�h�ٸ�&���]�I�� ��o.��4�����]�*�Lל�Â�l�Z�ť����1���̐Yz�y�~㹻g�-l����	��=�;�O�s8t9;���Dfa�z���}2kh�G������<\V�eQ%"�hf���d	ؙ�	��U����>�Qs�%�j�H��) ��V��DyO�̥�4b�fJjo�>秼1�0�
�JFu�7`�>����s��c>�����R��3��	��2tYs����UϽ8������N�S��R��w,�CH$��#�"A�L�s�����!]�G�YsUs,?��.�]�����߀��`ݶh������[�1m�T�!�N���r��BP�;�q��+�o2��Q�.��b����L��� p|�~fV��{3�]���/�ǂ�B�%�)t��'�p�ҡU��Ո�:��c\'�sb�8aKJ���(�Q&V��p�G ]�8%��ϒ��w���.��� �x���,B��(X�<=��O�{ֶ�C_͇.W'K��
�t���}_�p�����u	��suo���
�o��#���iMO��A�R��{��w<ۅ�莝�o2��ɕ�{�AQJD�m>f���~X���3Q��#W���8W{���m�B"��xX��GF��S��84���%�Y`�rts�aA)Ly�1U˸��l"Үt�5~�ݝ��uM�oe�׸���wH�_�LH0�{8宦�5濶'uP�����aKӀѐʈ��-�Mֱ-�o�h__���V�ɞI�P������m��Q����n�Q@k��O6�m�ѹ6�9��$�џh?\��v�#$6Ѽ�C�ݖ�,>�վ�Z�<���9�(�q����g8��^,��e[�\��f[�ۛ�g!;����Rŷ�3`��yT��E�Q�8S�z-��q"{��:f8�vf�i)ٖ��y3�f\v,�X���E�H��р�,]Hr���u�
d �GAĹ v�9�&�=��B�9�\�9o�}y	�/@c�ÛW�{�6�iy\�{$Y���=�3�6�\��Y�j����w���B&4-E�Q�O@�Y�Dd�0�[GPLWpVU��`d�Ra��!���vql�I�,[��q�&m�6y;^"Ǆ��=��m����x��Z���d�?��-�k�Z����ۣE(�\'٢
٧�݀ 6��?x�$H���z�߼�i�#s]���IH)_�	����R�7P�O�2��$�Y���:�+�})���0cK�*�"��rʖ߿1��j�Rl��o��hᛥ�1��[��I����^jh??������i�@��R���\I�c.!�����טPJؕr�<p�Ηi�_���0��J�wE����Ҩ����00�߇��3�>�#td^s�a�A<��t��$�6���f��w��P�G�s���%�{NLp���ʪ�̲�{�(B/dӿ�#�4�Q�&��bҏ7�n6>Y[A��Fg�K�6�$�!��
aN�����HϽJ�
n��PcKp����џ�u�Թ�� ��%R����4�VQ���v�=�S��L ��Ns���+�눵���s�-�[�(��,�6���g,��pj���~E5��:��2�����W�����
3�x�}ea��@��[F�,�u�Źc��,���+��H<�����R� ��lgӣ��g1��؉  .���$��dح����z�"a9�$L�c�t�/�!0�Č�hƜ�#X�#U��j���
�;�VC�׋�ⳛ$����7bύ�۽�[�D#o��~)�)=�B�+�x���S�~'��-���$+���ѕ��ȃ�J$�8��"�i��sd��~E�8q#[_;�W��u^��mKPs���ߦ:9���ߦ,�-�<�"k����[�@��'�`�Ig�F$��E��sJ[�$�
UĬԴb%���6O*����e.v�j3H-3��q�-Lw�y��Cb���K]
ԓ����F��E�Rz��Ӟ�ݯ�v�R>�z�>���'�~���g�o�/D�U�R@#�����a��g�u�Ӻ��V.�,B?��Բ����I���������:�;z�!A�'�1%<�����M�Y���������߫��׋='�d�����uE�(Σ��i�	�Juw�J� �˺x�*��C{T��%+�uq�wY�C����������$p7�4�hB܃����T��ؿh��*(E�ˬ ���(��E"�L��Z"ӷV��2�=���F�뜙ڷ�5�v�TZ9���p ��V���?hS5!?���g�͆��NcY�R0�����t��E�ȁ����,[���o�8P:(VDtц	'⌋eK����@;3�j��)TR������v9�24d�]uU�Hпe����NL�ޠ�v���x[�p*6���&Uk�*$���v��������DR
l���,<�t��#���6�ü���~@�'�`{*g{>���kn��B��7�+�d�&��V���bs�܎ͻ
��Ro�LY�t�-F	�F�d���H�Ev@0Q�Y��
��>ncM�����&i�&���V���ؠ���@����9ׇ�'��T�Eԉ�.,���T8���ӻ0�#3���mTV3T�|�K�@|5ӟJ��S�R�;sK��F.��;>z��ϘES�<[�s��6���w�k[��`ćl��0�ޔp�m<�R��M�o~oiP��0i�ص�A��K$�)$�~>�Q:65M�(:���
�|'m��\p�Z��.mm��A�4�b���Ǌ]�4mlr��0�`Or�~�}�
'�dQ�Iݒ�mw��I���`�q(�Se�Ŧd��Z�NQJq������F��4)�s�ȆS��8�Jw��R��0��y�z΁Z�[C"��{��N�7v�B?�}Kp�i��e�oߜ��gYB��k^�v���	!~祾�{�FS��؃̓�b��GU`|�jx7�i��QA�L%P޴rR����FVq�W]�~\4V��a/��-��Z��ݰ�]wmU}sY�£6s珑ll��%����c�?�;��mM��L���B|��O.��QE��3�y��4����lqy؏�Q�Z���� �'p8ʐE�r��`�Ɓ��x>���v���|+r_E�,_o�w�=����)>cVO�FZ��h�Cw2u(��@\߃"s�&���牢t�x�b���9F�v�?�3r��?w
��Y�k4�ZV�~���_ʒ�% oNs����fr����ÐX�t�����!¹��tU}rE�:��jR�Q�r����?D��a��F'�X�f��
˫1S�����z�A�O g[�g��W����Iv6C98i��F�6S��y���e��P.�yS���П>y��e�H�K�(XB�Ϝ�фG��X���C��F��0/���Aa��/���疵Av*��X1��qH$*%�t����O*�Qy��L`�F���1�C�?�Ŷ��g�t6���3�Ҏ5X1��@�;�f4�Lo�t���n�����**�@\m/cL�ߌr���xI��
�3��4�p�n azv��aO�͚7�-�'*�;^��_l��w�0q�p��
*�C]��f�o}S�+�)o|Wv� �	�q<(�ex����C��e~�ř��kUo��`�x���3�ð(Ի��]�B�8S��S	���2�#D#�0��`A�ۀ5���>��~5�G��]?�]9<^��>� �J	-uK;�P�ؤ��c��H�-V%�ꕀ�%�~,�����!��o�	=�)�&�{B�1}?��-���E��*�r�T�;T���m��T~�̮�p;Q��oD�(�S�+��?G��aC�/�Ē�yMu��E��1��%�? $`<]CD��r~-�cQ^��=��r��͈����$�}~�2t)�%m���Z,9)N3�W�sZ�F�O��0�7"�������l%�E9��Ή���J���\�����&��$K�����q����:�܆�ɑU����P�� �Bߊ�]�8�L�\�{��D��'".�7�������'k�|�:�v�q+e����l�Y�{Bn�x�=�9�G�R丩3�Y#T!m�x����ĺ�@����azk�2����:F? �[�W��bhhU���#�����H}ۯ����kW����p���RG��<+v�&ڼI2N�[�{�D����{������t5�"����1�-�jm�&�+�R�W(����_�VZm�v���ѷf��,�g���B����V�`��T^���n�8�)W��m����Lb�-%^�[VEz�>�S��.��ן��hS�OR������]��}�٩�q#lq��|��j��O�y9�x��o�~�y��~���`�ĵ�v`?Au�����sj�zk�dT�7=��.���3}V�n�[Ȧ�_���I8�����H*��4(�QY��5�cH�Ѱ��O��uJȹI��C,�c�BU�F4}�͘<�_m��!���`�
@f/q����	%{�AuW�w�,;�|0�)�h�7A�Z-�� ����}Q���8�>{rO�c�#�^�����]������D��̚�@�}�d����4b���-u"�Lv5��R�/:��7�G��q|	���|��6�%�p�SfC��#����wC�PtN�T�� ��B�0� �?���y����R��`w�ߴ/��}��ﰧ%��W�=�B5�5�	6�'��t�P�b�A4L��0|��e��e�W�\3.�u^�f�ľ�<��U����/�Ɲ��@�w��zu���p3���T�Mnl��Utۮ�.��="��<�"h�F���
'I5e*ƨJ�.[��v���ʰ�U� 3�nO����:,�']`�Oa�O�P�V�OL�56����ŋ���7fJl�O�m�~���c��_U���Z)���*��^~]@����#y���)�W[$������z�g�v�ή�4�i��v|m{D=s��H�Z%b�)*` Ҋop�&: u�,yb��)P�w8`�������*�u�������Ɍ3D@3�O#>���v¶6^ua��_h�3҂�v�GIc3ЖL��(#�E��!X�12/pj;"$]�B�>�M�����@ޗŸ��ـ�[���%Jzz���~������,�s�fϒ�g=*�t��݂���چgEύοT���F�]T"��W�6o�����n�B�	:�Q?xٜ�'���>�N��T���霌3?��1�:��n}�x��?�����������SC۞u�����)�'�ޘ�SM��Z���v�/ |��?h2�����@ο/�G,�������B�:x�̥ρ"����wu�;�����A�o�2Z�wk�x�ٟ?8�^*U��K!o�u�bt�nl�4��+�+�N�9�kX���w�������j��$�ٷ�+O4ga�(��0˩��%ωgF^_���·���Qs�p���1l�j{9��
��/Pu#
�=� x�@ʥ@�B�>�?d�J1T���A5:�/^���Uc.��/	f��z�@�	y��E����|��?��m$����*�io3G3y��O���c���@� ��F.f��^a�%E5��0����*4Y�ڭ�I�xY'�o�ON&1��(G"��9U��[�lP���PTe����}f�>�VXB��~��o��i(kP��3�MR:��;ġ��C�3�3��g9��^�KĈ��7��EFϤ�@�\h\�|]���)�b8vQd�ڞt����4�o�Þ�Y͓�
.Il�K���č��P�Z˶Z��g���{�G�mo�@!��A h�VDO�� ;�|�r����-�.����ʠ� �u<ZJ�i���Q
4]�������rӬt��i5#�[Z�&:�A��;-��M��,wu��� ���~�M.�ʿLy���%�7�Q��F���5i��f��(/O���*T�w�B�D�_)��L������{-̚2S�˄H+!ȡ��ڻ�0�S�#V'v�#�?#���Z�� l~��/�/�"&��j�����H'��?x�Խp��X>��4��"��G���9��N�Q�~���w���HBp���Q#��y�fv�=�3�,x���ț�:;\��;/܅��\�x�Y]ue_e��_IUm���j�+���e�{$�T���>=5��Ё@�^��u"�;�L�T�=��oeM>C��i?�I}p�b�i����ҡ��ȑ��6�K7A�H��6* ��۩��|��f�W��0-��8'gpF���r�XO�.A�aul��N8�X.8�t|���)q:���/�U,�9}��g͵̼����}��l#>?O���J����"��A��sgay,���c�vR�!���]�Td&}9
��J=��k�!7|e���in8�M"��__�&�FS��~����N��g�o�b�%����׫c���ƈ
l���{��1Ьyώ�--T�}�Ȟ�j�LA�?�~�4��^j_�Do8�*���yv�$�?A��;m���y+*=��3l���<|�V�E��IB�90���["���J�W� ���³�N9"N�>aB5���/5{	�O6w���T��]SwOx�ׂ�T}|剟C#��1��?iu�+�U�-����=4C�Ѳ���������I�66��䥮���`���k�H��lW���IBV��~�֮�'�M��ј&"_��ѩ:,L��NJ��<u.�E����7Vx��b:�:>�媋<��g��)���7Rrxh��V���GzH`�J=)���Bk{ҽ��j:�C&��pw�[&��"6_����#	��]�0�8_�\✄s���\���­�����G���K��*N(@#�B�;�|�2���͑��&�N/"��]\���iZ��ٸ��N�<}��pzb^E*/���7J;��$s�
`x���s%�Z�����q�Y0�1��-��m�Ρ�%<5«�_I%����~�.��Z��T���q:���UbdّhӸ��!��3+b��tQlW8�
�7a�T>u[C/�\ i=(�y��d�k}���������������o��� �eF�w���OH
�8�4�����G��~'T"���1�Ex��m:H��e9�9��Y����Ə1�l��G�X9��S�3{i*�нWơĽn-~ծ9s�Rn�2��_�
�n���re�]\E�羣
GxYG��9�d���Jn�����$�t���X��ޯ�~s9���2��V��Φ6(<���M��p)t0���ĉ[��1��� L�Y�D�g��t<�׮D���} j]�Qc�͸���d�@9/o� X�Ĵn����7��y���g9j`��Oǐ�M�vw��E���v�'��*�����y����a����`R�IS'��#�4���\�Yn��\X�㰁o��Z@&bd����Wx:�=&��O[�2']�H����N�>���7�:S}S/�v%r�f��֗@�֪��U#$.Ұ0.@QU�0|��/9���vx���Q�G����>t"�_̋xǪ^�t|vc�N��g��%�?&{8/Y�0`��o�~T�:c�w¢���X|���2�L��y)w���*���pbñ�S�,����H����趣��� �?%�L�N{p� ^W[�NsH=�I���6�o�O��/#}��>�'Bg���itm~�y��F�z3���+;�6�?f�	��7��6�ᇩ��uJ�r��RY�g�@�"����V#�H:�Ӗz�9���~�9����z�SJپg_��X��ߥ�R�_������-��1�NBۊ�ş�ҩ�MO
�$�g��wW�����9]��¿S�7/��t�e	<G6�� ������xflpå8q$�s���V2�8N��c��&s���]J��-Z��K�֮��a0��%yh4���J�K����HG�PvZ3�MU�!������}�ڊ�#��C�X�x�JY-0�	�U��H�V�,lDO����pQ��&̭�rf8х{o����V���N����~ �		������xR����X�Y�cE�-Թ�B��ވR���9!�8gbiR��FV�GfM�ݷ� q�u܎������A�W�xi��p�����LHX���w��Y����{ءǯ�;�x긳��^��ُ��9D�+�t~�`�G <ˆsU��T������/M6^J<�y��q+���Wb�5�#�����>"C4�冀^�a����5j��^ՆJ`�0�fB���D2�g-R��g�Q6Bn?���7�2-��ϗ��a9E
U]?D�!/i���\��p�:���K�Kۙ�^�z�#���J����f�\
����w�&̼7؃s��|�!$"��E�"��oe7<��£��f�]�	�K3A�%���$5�d2W���ç+��5����,�eF�`pO��B	a�ϝ�����DHM �NG���9��/P���6�����DkJ�2��h��A��&��aɐ����u K+f}F��|{lQ�|����=A��ɐ>q�؇n��+~�^���l)�vjI7 dՐ�b��gF�����)�<��a�#q�f�f�N `�Q��.���1����Y�'�˚�Ǭ�-�!&�gWqo�F�!�X[�m�%N>��#2"�6v���8���T{ⷎh([�9;�k��˕b���gh|F����4�q�� �&����`�>��3�tB$����^�wDq<�%�Z�8��{�D�z&�hR�I������� �{
����A�I�5�'���#j��i�J��fx���_�9�@��i=q�gPԪ�g1x��{Q˓����~��ҫ��_�/ZF��E���j����C|M#W��#Z��M�����v�zm,���-u���h�\�}V�Y���H�f��[2�-��Ac�$twKCc@)8k~�'�_�����//Ş�J��qmҫ��7���F��.i}�0�M��B��.)��Qa|>bd}�W�R�?�%��#�4�\u���r����}��X�Hɕ��Ď���F�Yp.�e:��Y��h.Ry��h&W%��qM���CjR?��4�8!A'���z�_0%Y�MV���q���C���e��8�#H e��U�������2>�.���/{�����'=ٷM�3��
rV1�W����6Y둎dj=`���P�O{�*V���I��Mf����K���ེ���!Bj�K.p��i���1�� ��Q�q���R �5���-���)�vَ�~��5��h�-/k{��V{�������I�P=ƭ�S��ƕ(0���)��,!b��q��G �1������O�2��G�V�p���4;�)|�Z�LF�쫮�{�Tu��O��X��|�s�M���F��
���N���?<(��9�[t��)�(m� 7!����x~v�Q��J�i�	���Co���$�ȇ��c���'*II�/4�ط���a�*��j�0^��
�1
�vN�ҫ�v����^�4�\"�y�<���8�9�r�d�E=������=���E��k�L��J5.�I����;R�*�p����b"$�^QrZ�#��RPh�~���pr�}��=���������=5�O���0~���Z����������ܽ�i}���,[ ��TّLލV{)c�(l��X�m(������t���{:&�t K����RC �i.�a��ZX���j��'�����,|�:^S��9+l�)�ͼ���lv2q�<��	^�������,�'�^��i#��i��=IC������ΰ�B�0��V��~�m����p�ʚ�t�(���/�h���A_?e� Hz�1����6��V�V�Ξ^�D���J8c���`�Y�y����Z�o�(EL!z�&��%v8M���|��r�Ҩ�5(�F���rǁ��X榦��wr�5C�Ta/3�0�� ��q5�2��l?����T|�2vt�D��չQ��8Ƚ��Cn�*jS����J�b4���kvGk;�\����M��1�MN���
���`O�Bgx � nI�5�y���t:���Z̪�;�qnu���	_���:ED�y�6�m|��\�^X��h*���}hf�6Njh��>!3$y�2����Z�����͂�omS(n�EJ��K��蝀="_$���h�ӿ4�q+��Z�i�8���K���܉�v�\��Ba�;�[���$����	F��
^�%���AӜg�t����q��`�в�{�&'#ŹՏ|��P�щ�p��m/�33����7�~t�,�Lf����~�ڮY����l�������o���~�89S�5�u <��Q�-leB:��h"V��A3ǁ���>[���"~T��U���:� ��������BDi�A�Ŷ 7��������pU�����x=�_�rmw�R5-�[
�2�W\BȉIa�1�Z���W�;��@n@��5v�~����zW?p�q#�X�L�F��
K!�;��Ĉ,	��3gv(Fxs����s*�|�������'e#�t������y�8E쏳�,�27/�v��{��싽�k}�%&����ޑ����Ӳ�lH���exL1`��M����)t�{K�/rǛ��W/���N�?a��+�/8$N����sS�c�A\�a�Bڗ�S4�'�?R�����V4�����Y� ��ã_`P�F�{���b�M����@,c�� �b�J�}�YM�)0��BSB�݆�J�$*4�9�.� �L%���~Έ�h�c�[G?��g��T���8�F�fJV��I�]m��D��DWsZ\��SJ	l,��� �u�TG��<�`���J%�I(�:1pt���e�w��j'���Th�G��9�]��=&W!;��i���k���=���r�<4�jN.��bל2�VP�	
*�צ�=Y�:zJ���ȫ��8�*��e�������-��^�C��/7�ʣ����j��������~�"��i`��$`�����l�%���%��r)́ G3��K�w!$�4*��/
�r�{�X��_�X�-�c��.W�ݖ��e���}�w(�t��^̰�������`�-mE���$=�x(-���'��U)ۚ��[�mL
�%��@Ĝp��ݕŹyϰ�����)DnM�c�9�]Q8F���U�g��*1��ǧ�E�#DI�	oB�Ѩ��t�K�2��A
�Q��)�f$B��`��S�p\�%,�4�4J���7�x�`��5�g \x���6&��r��M>�t�Q�U=Iwd�j����B�����"�VyA��\���.�Cl����*U���<�UvQl����� �V��x"bD�gL����(S��5�Φ
 R��	_+�޶������S���t�^%�Ȫט�We�ȿ�i5�O�c#oZ�Q_g���w|B���e��bI��F:�[�(��@!|�L���h�ǳ��	(�6r" ,�bjE����B��%&N��ԏ$��d��'��[��+�[5)����)� ~O}U�XT{^C>@-�z����P��h���{B���T�/��II��u�`���xD�0��Si���kL��?�kXc�b"��T�A�fC����mDoMR^��d���(������qT�&@vy8h��|y�w}�W��d]Ƨir�N��6�������7F+H�*x"C�~q6lư���?<�cvM��諈�ͪ�b��Q��WKVo<Qz;䋯Ji�S1+��9c+��rݫőkV�Z�.W��x��|�r����>���j��\�j!�	��^/&�2�yXV�ꃲ֫�����3����/�1 b>�l*T�#���Ye�(��g	�F;o�9��j�oj���� �󁂈��b+��KL�Ր� 7���eQ��Klg���لP'+��������N+��K��M�W��b��R^�v����ź�uv����f�nA8(y]u�䕇~C�;�#/:S=<hn��n˓�D 
~��d&H|�q5r$�Ѭ�9�h�/��8�K>����\�鿳%=&��BZ��,�=R��9����6�ZK�Y)kۉ��%CL�"�O�;:Jm>�Z��Z9������3d���P��d��$x�qq+U�ǧ{-k��}���J�[��8UTc�!���I���j$�<]�"���S��w�gp��1�
`��p��Oߧ����T� �� $�%���G2OF/����X_a{N���e�2zr���>��O�R)Q&�x���a8��}˙� $�.K��]���ϰK�Wыp�]�]�$g��$�bfgH�/.�b^�
�f�j	��U����_B[��k���/�k��p�i&bg2��a�^q��RMl�aգ}�h{x��\!�[E�ѻ��@j��۔-�d��ĆA�t�<ȥ�����R�d���U螈����#X6/ù�����|�B���`��@ԠC&欏��������
ɟ��$o�P|��ڠ��y�	�u�����B+tD��y|���6s�߄������C��g:u�RG�t���ʶj7���睚l2dE>Ix�d�3lS��ʂ���*��b\{,�^~���d�B�������W��D.	B�T%g�7QJ��� �&hb��=��k�)]�]��fF�b2k�`�ip"�)�j6S��P%,��m:*�c�~���T�o �R3,{��e�j���-����̘:�k��	�=v��;3�
��T�/�����tL�W}o Ԅ�Ů�X��K���M'S��R2�-�:	4�7�z�A����г���2�p��%�q�
&��Y��`�;� ��=�3c�Dp�hi����e���]����W��,XV�<�������S\�h�Ƀ�:�k�~qT<Y:�~(�*��Ԋc<$7��%�����Y]J��p���#��噚,���^_
�%)���i��+9��m����$��Z���\��!sYQi�e��AY] �8��ph5!��f����k�툠^�n*p��o""� �?$�K {7������Uq4v���SQ8����"�9�
��4������=Y�q��sUo~���i��c��	���3!�t(�2K��m�#�Z���������ʘ�p�\l@�S��F�f��7�������OM��p��3jK�X+M�qdc��!dd�� s�v��>h���M�и?B��n��H��8�On������*�@��:�	�� ���D�U��^�
O7׳����l���iԁ)G�ߎ~	��Y�Ϩ�G%(x�ґqD �,3.Q1��@t~A�8�
�BƘЦbW71�9���9�KO�oV����03�,fnw��tpP�2�m�J�
q�LOC��q߰�/�(�����ϕ�Q�9����%�'�r��Mk~���B�F��0c�z�*��C�n��'�y�R1v�<���g�ɞ-�� +�[>��q[���/
�w H�P�����l�9��YP�RX(a2}1�7b'�*�ܐ�� �(��H
$����c�(����Ӊ	���-7��=�X���M��B�������qg�G�MG�h�M	��t�_}�%o�K�&�@�ǩ���3D�/`}}���9�k�E���F2� jI6���
CM^t��� ���>��:�������`N?��L�I>�e�b�Js,E�iOE��,��P���y,�\�>%��4�RL�?���V��עӅ��f-?��a�2U��3/!��?k�@���*xˬ�)���K��7���v�2��5v;�(fF�O�o��������1G��{�#/ZE�|�d/��dR{n��`��B-+�խ��~����˥�I9��N[J�s�Z7{�S<�;"�p�
\=)��U�H�����"��7[p�R�~-&!�&|��9�(f�������N�`{)����`ʋ��F�0�Q]cY�x[� ����Z���3h��x`�����WH�U�};[Y)����nxݍ�RVn!�Z�i����(d.����X�m'q��a $�3l��������A����%�������H?�vW~0Z>��SFԳ)��t����p�U �8�;�ɖ�D����3nv �Wc�A�pB���5tI���́���Ds�7�w4q;�3��Y�kW���\<�� )���cuP��$�ؤ�ϩ��*�(�5�Q"��ؔ���R��
����qb��'ȮG�r7N9����B�1|^%�o�S);
�KvDr�~�L	r�w�PzH�jqZ`aV�܆�C<W!=��9bQ˟#��M�~K������.Ҧ<z����"o%pv��]��zDR�����䪐b�Pg�u�����n\�'��w��z�N�\(d�`���<>�ѣ��[�4,
H�d-�/��{.��RO<dX��� I�T��ńĉ��:FYJ� Z`�?�ᘀ���VّO�r�Hӧ밿v���x\=O�](Y��99�G��-�[easeX �q��կB1)� ��������br_1�C��B��$C$P?4�V��H:��0��u�"�v�uݩ�f���N����c!ؾ��AM<h��bKDU\b�A�YI�--8r���!�d�=\�v;xry)Y�M7��x�x���U6����K�Mx-��o���Y���oM����YU�,��L��j�Z
^v��Px��װ� �P2�>!N;�yƕ��F�h��Yz�##��X�q�8�;�?6�}�L��ļ?�ho	�ɳ�vu���KQ�
�m���Sf���3��lυ��&Y֫v���tL�\[�����8���$���2,!)�w�a��rÔ�0^4�HQ8�|�;�c8��8r��V�0Tl�C\Л�Ŝ�X�������c�+�fV/o� �4�������{!qn�*�ɧ�[�%����"LZ$�z�D;C�$�z}�u�d�Cv��@O�|�r�O>�H��x���zY<��cs���﵌Ri`M�8�O� ���ͭ��,5�4��H-A�x�T���b��g�#�V��#R�� ]+eKZ�5;O���g�`�b�*�7=�F:Č�Yz)���]Y�n5�鐆�[�/ׇ8//�~ģ�S� _'�����:k�@�w��P��!�0Dx�b���_�� ���m�']3C`'t�{�J��H��/- �e�ux���+[����:S'���N�j5��T����T��ț6fF�
�[�H����WW��b�˪����jJo���
�_t�n<��(z����R��S+�Q8�¯���*��� �pD�����ŝ�\�!�֭�թt��*O��猐y�A ���*IA$ɐ8����
㕭�j����?>9Z�H�8W�S)9�o�d�%En���@K_>��d�oN�u�l� B�2:��������C��+����P�&@!�'ӱ�w"�Ss��ܫ����Y.G�5���I�A�闆DV�5�`7�y�z��-X���NX�GU嶵�|fĮ�w������ʬ"���\�}�ݽ����\�@�M����7�����y=Z���i\}	-�T���)�R�(���μ5ꯉj�1Tf��3z�ܨ
�W����u���� t1�B4���N=&Y��<l�K7=W��>�F�A�À�*I��l+Գ�m4y��}���#"i	�����3Ȗ�dɇG*E��f{]�n?���T_����_ #�ujudkZ�����-s!JER��%
Ԛc�Ԩ�q��U/LWpZ���ǜ\���"��c��(�O�W:�!�3X��>������^=�B�AEɱY�#���vb��J^��TA.�`|L.b�p(�}ݹ6Ӎ#�L��eP���(hyd�9��%�\�꺂-[�T���o��,$���+�u�=cb��G:%��+�G����@DƁܝ�_����_�쁮A�?yүbN{ȼJOΩ�]�}�r������BC���f	I�_�/M����0����*�E�Mv-�s�5�WR�1��el���k5E�D�0�/�7��iD,n������SW;��췐s?��k����̲MZ�&��)۾��),�����֛��^��r���ˡ}�mYimQo��t��F�C~l|m�^���U�=���B�����=��b��1�"�R��>HF ^;�� ��1�����KmJ�az;j�3�����1f�#���V�Qk����fΊ<�M�a��5N���7^�.���U�h�V��үy�+�Iu���$`;d��"9�:����b{i�K���|�����˃���C<�K��7�8S.��;����
��Q��7C�`��3�ڮ��A�Uv̝�o��M�X%T��l���)&� �e�2�lsr�n㒄��}�'��N	�y8�/��q1� 4�ʜ9F�l]1U�}Mn�O�S�ritt�������7X#6q�����i�"�L�3$�lGq�$��c���W��A�֠����:�#E��jwI3B>���,��1��`Y:�2HK�~觟�c�3��X@�.�W����a��bl����k%i��-G<�]��)|-�(���.�~LD��l�c
O�0c�,����1�.+� �O|,ڕ㲁XM|����j�ͧg�����j�-�V@$R�?�3�e-y#��.\O�Q�;�>l[�U�Y��Uδ����粮��x±�	��z�qIַM���9��:��x�_�p��Q��!F�E�a��M껁�]�l>�Q+�p&B-E'�����J�sb���1V)�C��P	1((��u��G3�1�:�A@!�c��K4�g~g�MK1��B�_�ez�l/����Kִ��C�u&��[෾���o�Gp�v<��^J�߉�5�Ó��$Gn�=��s��T~jE�vP�V# �e�"Ͽo���fR��
�����@����>��¤+C�g-/ˣcg|�!)* �����hv�,s]�f'~*T�=ǃ����|y�"�$㞖��aظ| ��GK�ˋŉ�߷6�ޯrQV�M�A��r�� �miL�=GXJW&b
Ԃ��A�������xŹ`�٣d���a*�=���3�]�{!��J{,TW��C��Z�J�z�W42d��{���
yaj������U6.���$�.cy�0
4�y��u�nͬ�i�1�mKu)��:V�cl���)"�����D�m�ռ@��<�cG�7	����7�fr�_A�A�R!!�Q:�G���\�e���Hb��d+e1��%�v�2u�(.��xF:�h%S�9�*"ވi���R���d�F:,��o2�� 0_i���9h�mw���N�ac�����p�j��pm�@�NRXx���V������/ЕT�o>�~�"�Z�%b���1��ȴ���	�w�0c�]@�|!�q��CI~�ѐ�?�X��Dߟ��<3m�Z�s��n���)��ؔ�i�v�ó����,��,��� A<�ơ��qV��69c��ߥ�<�=��6�;n�l|2n?��2}�/Ɨ���=�������rmo_�j_z��RVf #�Yv�o� ��Sj����A8��W��.ۥ�I�~W���Y����A9n�TJ���x:�Ò�'��n�@3l�1 ���!GZ�+\�7�$����I/�_�'�o�;����O/�:�o�Qa_�@A(:\�������e�5���b��ǒXV) ��H��O��`9#,��x잞��Y����S�f?r=�B7>��b��W�n�����d8sL�e�[�j�]S�p������#�z:֌�[~�J���Q](*w�W"�9T�TJ�\�zK�S['�GI]&
@	��l��{�a+z`���9m���Lq���C����F��?���M��E3��U�:�^�Tu]m�"`�qq=IAQ��8�����3��*��=��SIv'Thlma�� �����"vL� rސ�H�����g�t�?tͦ-�f��Ra��i��<I}^�2�DU���B��(eES��>[�*��S����=9��Kl��?(��*:�(\U���jJ�T�
L{�K�A�&2���}eΙ�]ɪ�y8��W2;`�Ioz�;��`�I,8&��{խl�N���t�L��𯵉��(Y|�z'��=��Q��#�;1<@x45^�PF�w�LH��a��2t��?Å������B4N%��jP�~�n<��9�٦��AWV�=ÙL�\�u�2��hB�c4����D�y��GfSȞ`�f��A�l�2�Z
�8|�3D�͊1y1��r�XQ>Y��C�#����xHQǇ��ڦ8�+V��:��DŻ�b˸P]�bV�j�w��`�k`z<!�d=�O��k�����]�Sx^�!��o�H�#���zO�!�� О�u��v���lj�m�
�A@��x�X�m�&�5%3��E�֌0���~7��4:��h�0�7�^���7��w��R'�9�����+b�͒'����x�O"&��~&���uj���K4��@������� ��9�4�H��j��4��33Λ�~C�qJ.�����x�e�Ս�j��<���WL��e;|B�q;��G���Č������|��P?c�G/Բ��V\�*�X*Ǟ�sT7�rMj��� h�U�9	�V�X�=��u���6��!χ
�,|NjR�Ŷ�*�M,?x�՛�-
Dh�l�5�Ӽӆ��^fX�ǱR�8r|�l*�`X�I�Fz9"Xq2��Hٕ�]�L��'��9��s�J���7#�]{��%�p:c�6z�^i�B�M-b[�!�]�����CU�<�k�V�a�؁1�<i���34��ߜ���}��i䮈��:R���&ɔr�E%�c��މ�6>H�ޮ�"��Q�`����5�/B')���yp�ch�a����������%��A(����٬}}|�v ��}"� 8vF֧5
�j�̑�V�\�AW�=�  )@!x�ڿ�<w[�:p��K�u��z9�|휱/s�9�^4��s]NֳEՕ�'�H��zQ��p9��Lʋg���?d��vk���>���*\p��#�(�(��&(M^���SB�=���]ؔ7=_����xٛkgԱT��ڼA =�ج��]R�Dh��q�yZ4?n��6H7UY����L�"�a뉟! �&_S1w�TjL�5✄��h���o)��ͼbiêY�k;�x��G�(I\�[�X�@�`�`\��]F�s.��^I�꛼�I��Ԯ���͡vl��[u���\��v���S�+�w4GxВe}��w�y�1_�M퐗2�bw[[6�-Ec�)?�]O�۸߳0�K��hd�JM�$�1�A� w ��'Vۥ3�s�]kh��SZ��Tqϕ<��a�	��R����՛�x���4�C���	K��-�<�İQ�d&���Tt�
@�yڲ@P�lFt�u�'tC��t�X'���bh���9�o��\�"���7�x�67�iJd�5���WŘ���߃�Z�db%& �r0�8q����eΎ^�ю���b�3�w3ɪ|h�p%�Eo�onR<��쏈����3:�A�'U\�yP�'���%8F�Օ ��7��Klo]��6����6c���<x��:g�4��C���Z��1���te*x��v�E�gU������H"��	��[�O�_Ws%�����LyMm���������j��'p���+<��o��;�P�Ls��� ��Lu�(�V�k���`���c�I����[�	us��'pW��o��x�~��M�Piоj�� I�E�.┢�V��f�Da�M����tu��q�
��3)sx��u�n1��;�Ϡa��q�I�
 �s���az!��Z��e��n���������H�@���,L��YqC�]�~:��tޜ�n �B���yP+���Ʊ��.?pƃ(]��9�zbI)muR�s��wM
+!�Rls��TҞ����t��ƴ�����I��}��g�����`Jj����{	�c6Űʶ � ��t���GF%�8/����`�A\��荒:��I�3�q�� �v��%�c�D/S$-���,A}l��l!�lUO	��A�,!���E�Q�a��@1V���l����A��0��X�V5y��=j��!g�if^1(��7���Z��:�-��Or�A��??35|�f��c�u���8�:�����6D+�O�,�;�Voy�`�#�&ёj0Z/�\GA�4��CQ��9��sl��Lt�Cg}_i��#e{�H��yKE���<�D�T�P�/|�>(����,1���1(���o'"1&�AD)�CM��x������Tm�y9�*r��jQ*i������ܹ4B�VL�;�L,���[Kgq&������7�kР��E����®�k�����A�/p�˲�G|�N&]��,3	St}��N�Vg9#>O<�ƈk�D�����D��w'��_ރ���t�y�h��Dt�=�_�i-��R�/��f8S�f*�2w�d�E�Bb���N�B��<�����E��Q���k�a�S���� ��s_"1?b��h/iN�Ke�J� ɢ"UN���.ۑ������yQ���1�����k�"��������g����q��o�ۻ�1P���:ѹMp<�#�F06����z�|�R���ʥ���s=h8v�X���}��Jhu"8�=)K[O��W�W��(�R�ua���;�]�28��4/N'E}��/}�v"��d�⡆D���`G�}Xb�ZO���|;
�]�y1��u+�;?�g���2_v	QI/�<�,�*^��������D���?<�q��b)�a;����p��έCO��M�e�@�c����X�Oa�K�t�����>����G�����o�x�����$ޠ�$�$P��� 8ܦ6������]=!&=��� E1��R�>q���um���ɦ���t�	}t��[�I�+F���3aa�@D�'lF�P�0AD ���3v��^�:U�V>,B��<(4�h����0�38 �,���~Y�m8r�rh�ϝkUl�bvL+$��p�5����<<h=C�$5lg�S�4-����cvˊ��7��@.��w�k�����T�2�虙���"I��)2��n�M�@�9|�u���{w��m���F}�@�c�g1���a��"���n�Q���:�t�֜�r����?sXvC'��v��axI���:�N$Z��CnX�ĸ�Ľq?�WA�(����r���ӥ}��߁R�	t"4��'�r=0�kW��DZ p�`V���i+��4���"��R�梙��ϒ��H�߆�>������<P�d����
{>Z�NW���/W�I���N���|t��{/�F>�}n�q�0���ż <y�f��֠k34|Cɵ�R��ת��g�Z5�u<7��.��ι���:�q	V،ͩ�|��esG)�k�p@�9X��96�{� ��+|W�������LlӸ��A�4��	��|wi�����v-�Y�0�r����X	u"�K�qo�2$e��<D��\��F��?���Bn�"�[�FǾo��9觪�2O�|/����$)^�Ʌ�8)A��V��������m� 1��O(�ѳ��D�=?��ǒ�E�����j%�>�_��(�ovm2o3I��4�x��3>�?;Ir�Ϩo4�g��a�㠎��u��<v�p�x�@���P��5��s<�§gj���Iй�r&_��׾7X�>�1-���fp=bNr��qw�A7T��N�jgS�^D�N��N���Z��-���à�;���9��pH��XkNdU%�k���-d%��>�_[s>Ƅ���7,4s4|�I�f��<��8�NS�_�+���y�HL��)1X:��j��a�5�@t^sG� 
\�]"��be�o������ە,ʗ7�ݖ�c3�� �x�#��D{5��HNL7�v�]p:��w��.�_�����@��f:3\�G�P�ơ������4N\[�H�>z��v,�:W)�]&_-�E�øw�܃r:;��d�[���P"�J�탖IZUXZby��(��"�fiBY�y��+~S�p�:�К����{�o����f�����n�pGi�N�y�_X�$d��q#]#ڙel��X<<ێVl"٣�����r��9�ѓ�BB�%��3��Jc|!�KQ��A��u��Bj4#�/�r`��i�c�����~�f���m��oF�+��(ݱ��~���!��e.H�R��*�2�'��m������9b��L� ��U{	�����%Ҙ)�[����q�m���,JXRJu���DZ�� �6"̽�ciCw d,K�T���6�Z
��L��{L=_z�����w���><��U��,�
�L�+����%٭x֦o��X�-f4N������
�	\6�<��N'�WW2�#�D��v�����58d�����"v��BU��(�h[�"La$�)$M������l�|�̿�=b����O��Zeu�z�'�gK
p��5.�W�입��!:��O��~��pc.Wv� ���]-@��W���l�>����ض�1o[�(���%R��&G��=� �P��s˔?J�j�*�$ �+u}'ZcYY����q>8BQ��F�Ya+��3g[��!� �9�Y�(�}=�ͿA��臭����D��v^��]<
e����_9��o�Ƞ�T��š���&�2�a[QxG�μ��Z�wx�"�BP��u��UbF�ֺ�M;"�S�D��v}u�7��Y�pф#!�1��U�pXV��������Fc�uܚ����΍C!�����1�@$U�m�6�gM���PvZ�߬A6:���,��4˙}J� J�}��P��m�r:k}oX��6��ͧͪ�
�ﮖlu�=1\k�E�^���:��[0�/��s�+o%����|�)���d���)_���[>s�p����Ft�-�����dؿ,Mz,��^����Q�.Diۊ&���{��w����]��k�� �u�l�Gq�����8.�c�}������$��~1LR��g1���R�%%6Zrѹ\�-z)��W״>�SWi�dx!���3p�36(cb�x�~\��]��?�Œ�ā������������{�Puߘ��Db�ǟm�p淇.�b�3ۮ+g}|-�^�c}A�P�E��&�n%�猬�������-���
T��j�pE���Q����*��/��u;�O��v����pDd
,p���E��繸����80L�`�^�l�C8����F��/��]��!�JE��>�h�\]}}3�JxZQ�˛p�akn�6Ys;���EՁ�h���o75$�W�5v���پ�Ǖ�. y&˛�`Ǳ^�r=�s�rQ�1w{������_�����އ�<sȆձ��a�@����r�m��Ȩé��4�X��� �J��<z|�̮�&ZW�
	^���b�N/ӥ>���u�o��5��gYu�����+A�)b�����-AIG��@?p�0N;~��T�
7O����,J�C��'�p��Ɯ�i�W;QQ��@�b69}��"' !L�P����]i_�u��e�$�����O˗��b��"G۸i�+l���ۮk;M`�Ѽ�VG/u�-s�S�a�j7D��{m�FC����㮢/�u�a�n�ʦ���+g��:�0�f�̌�R�wԑ�����N̑���.rD~�5�X�3�������F~��7|n.7������ɣ6�
j[��fe�_���8�X�����/F�x�����X�0|(��攃�:є<���qu	�w�q2������'b\�U��We����]�O��O,�nL��������D�ac�����H/�_�r�W YoN�U�D�c��5����wa��	J��и�5��%PmN�Xs��</YΕ	�J���̎y�����g�jU�;W�	tY�(�kսk��K�܏�����g�ׄ�o�;^#���a[����u��|}�^W���s	<bN+ōkm�HE�m��f&��[�,��V�=�[F�m�����Y���{cA���v'��g8dk��5�W����|�_�Z+V��X%�&�S�����ƷՊ.eHUZ~vO�l��Fa@`��X�[�ߴ���h���� N�]0�Q��t�Ǽ��8�1a$��s���g�0-(��6�?�껱:J^�i�ݴ���;��V~�#!gͪ/���b��~OBmU��/XZ���lOq&��X�B��p F/����_�,���/Y&�n��;��E�)���s�Go����A���������jN9��e�6|`կ�����o�G؋�F�q��t@�IU�-%��_]=��q�.�!����=��!d6,"�NT�g�Q�#���A�r+<��[x��s���X� R��C��/sc�W\��=�8.^U�6�\=���]�1b8P[�
4lV�_��Ϧ�U�*4�C�1����f.Q5H�!��oϜ���O�@t�[l"���ԿIP�����Z�2��%���ᾂC'�}Z�����s0�dFpx2R��NB�`S�y���-tN�q��E��ZM�(�7���	B�'3�m��aK~��!�\"�"��]�Ħ*RO6D��|{�.8�*w,�5�=[ĠT�y��޵"�͎1?E2 ��}P�&"����O���$��R��<X��aͮ�8�l���]���v2s<��D����C�S��*ih��'����{�b�I`W��W9du �����!M��>$�Zh�<$�ܢK�m�X�C�JD`bLw��� �|��к���Nڊ��̂�@*6�|%Ћ�LH���b�S|�$�J�&�+�h��˕�}�.��5A3��m�<B�.n.��j\e=&�Yg$�n��^,�z.�כE�F�)�Rr��4�u�w.kaUz9,U*��L��*Am$7�A�P�^��Ϡ~C�z������$�<�HF�`$I4kz�� rs�i>oѸ *���#��<m�/����la0YS-�R��\(;B8+���>����T�AS�+�(�.�tm�ɡc�̺t�[I���w���㔼���b��0�::�<t1+�-��C�HV�G(�f�� ���v��J�	��Nq�m���*�=\��� ���)X�`4�{�tc;'}��v��D�Y�7N��6��-4��g@����+�\�B
�G����ZY ��R�'?�I�N_�l�nA�(?��3n-��˯��F�*3oّ��Ͳ�Aʫ�$��`�v�
rEg���<�g�۔��K��r��W��顢/��/�C��ʕ����;�1p���+]aA4��@ ?�6%�b�h!}��3ų���ɂ��p�'W_��� GQ�������ԫ"uYQQ��ݒ�+�[0��'���D,�ܣ�'ԚPRA���@���"�9%=��y�Â_K)�I�P��7Q\g��C�6�.�(�YSk����ܼ��Y_�$���V�A@ٯQ�T�E�<^c66�0��s.+�j�^��:ea�3z����_Jr�/r���P���bSشp|����ZY�����<��9��CBn�G��%�ۈ�^.mK��k��C*��GA��0r�,謎�o*=L�!�P�H߽�D'A1�z��mI�C����0AG|�C���6���& {TO��m���r)K���L칪yݶ�R0��|���t���i�I���+�.����$��;6�gd�|�̟Z�ߪRZ*H;�e�.-��Ng� %��~[�{Ě�k=o�ac�����?q�|��><;��kуgN�"��,����wF`�8����s
���~	l�
Z9T 5AYTť����@h�����AOU��pI-��Q��z�7�3{+�T��s͐ʄ��Sܞ_�Y��,=c�N��O@]{�8�(��!�h����6.���>�J�Z��o�@�XV�
?����?�j�y�k*Mt���^�*�/�wGg���������/�a�5"�f��0��PGT��!�����6�[t�{c�'`�H�`�֍M�M&�;~�&Ƽb-~�4��b�_b'T��D��Ĥ��`o�@��к"�M3=��ى��_�|��u�ԹT�Jy�g4з�k��7y��j�v4�jӢ�5�J�8ȭ� ��m ��L��7�����.^�zѣ1��}We��UK4-�@�mj�+��B/�mbJ绪��#�"�l�w�K�|?CPK����3��N���˘P��Aq*z~��j���R �'���-��!230���_aa��E �����)�z!`�bFl�����3��pY���ܡ�u�(�A�d"�PU��Q8ϬT�: e�rjT�^p���ng�'jް֨[�Z����O��;�46�p4i���nW��S�w�����TДC�X�UT��9�fl�S딠��$$XTtD��և��s֡�CKz4��4b2�#7�v��� �A���@�{�Z��Q�xU�z_9�F���A���{X!B[꽣�{�Q�b��!-�C�{U��6T�g;tnN?�yU���l1o�6 ��D�eia��#��A:	Vgz�#׻N1�j�Rj4V;֚���K��R���lgp�/�⥴��U�w����M��]��'H{��h0��j!�i�D��b0r��hJ��=s�=5��
�A����_����2���s ���	�L�9��qÆ� �f�$�[���=�RR5�D)ݝF�@�s���6�����+�O�*����XN�ܡƀZϦn1 & <�޾�����8�O[鼗�y�q���KcI�����-�.J�t:ʜ�Vq5PNi�GD���ʲ��ہY�(/H��ZA�ǽ�wA��N[И���R0�����Z��58�C3#ߕ~R�{@����ՠ�r���0R��09דhg��(7x�L�	�Ω�ă�����]����?�aO|�ʻ8�������`�;a�:��.T�[�i&�ƒ3"����]N����P)*m���,��H���x�
BK����Z'�eR��{�zH���P�a�Mh��H�#�+y\��O���p�������]yv�U�Ao�0�K �uv|�� �N�j�,�e�p~H�J`�w�.$-�>7�Knt�y`Q� ���s���C��(���DƗ�o��^�
���۔bԾ륿��*��6|.GQ9?���M��
,�5߯D�fId� �v_[���s�?�(���Dq �x{|M���&�!�����&������9�4r�*��`ͤ4�ܨr�4e@�Wg2$f[�qE|�L̦�����m���3�=��jf�ŚT��b�{��V��Q�2ōLez|�4UD�ʲ�Y��ߤq`r�U���*P���$'�]��d��q��S�>^�IPIq�����ד��!��v�s��|����oA2�s���)bqF������ݍm?�U�,(�A�z5J���G����������PF"EA�rWS�[�o��hS�i��*A �PO����R��)��h}	|W|�T��R��$Mį�`�=;��b��u�=e&D+�&���7��3�C�<	�$�����0��*����!B{�$W%�ow�1x�/ ��{�;�3@���@Q�!}p�EA��T��%�}Kq�2Nmr��e��PxU���
a�a��K*|>I�i+�`�����ĥt�6v����_p~���kx���Xo�|bh�c���2�G��H�6�R'�y�Ϙ@'�uWh�QJy�B�����1�RN+��!Ҟ�w����"��h���;��,L\s��:~����kϫ�6S)�:a��'_����Sl��9}i��"wY��a��3%O��*w]��u�� �Jiׄ��~Z(���?����,������J�į�����8�m�Sĥ�N&�ʨWbʷ���/��8:ޕu�C`8����C��G	]yF# Q1�����rO1��z*�
u~V��M�Ud�4�B����<�F��7��4!y�����=Mj5/�U��_� ]7iZ�������O��4��"J�fn���nu�	�M�-��}/ gz 卝y�P@Tq?�I���!����� * ��;EjV���a���/��ς�I�!g2&���&���[�޻
�Nɩ��ŘA�����c����-��J�\�[�K[�����.�j7z�&�G*��n���K�|�OAm�/�=�3�u�3e��r4gI@�)E/ ��!H4����6K7uk��m���(�W�� \G�Fh�˙�ؕ����Y#c1jCV���2D�]Ohy��)���ϕ�` ����+�ڛ#!X\Z��4^˃Nj��)X�%�.�z�X�����}y�=�9%X��W�	��c�aFې��ǎ� �~�!�Qf�IwoH�e��")��z���������=�i��$��/�/���6�������0���F񯧇:(����-'�e�����dĭD�v͢�-Î��L���l�)�v؝[.���^���HA�,.Eb�s��~[z��4����k�J��m ���h��~`$�a�h��]�T�`D��H��2B�a�_����ڶ��=��>�X~N���ju�*�V&̦u�ě�� �g�����r�A�'�/�3=�R���K�DT�)���'���R)�u^B��W�
�x�aq��Hhn�� �}��痹6'�.Xo����o��T&�����LG��pR�n+@�]�G���X�x\�B��
q �r�<�������A��9��mM-�0
Rs�".��@l��N8�j�����,�G�k(���j��;��x�9�i�1�K.�iaź+7d���P��y�ƌ�Z�b0{\p^y	n�FĐ۸� X<|�3)i�.��/�}��a�a9}"�N������$�{Uj��B�c>��$eܾ�NO����#��Q��4�ԧܙ��ԧD�� %-E�\$ ڀC�#��d�?�0}p���7qN�Kڐ"���֮')�$�u<T
]*G�>��¼�z�;��)N��T	⣬��]�<�����B��|D7H��n�G>[�k���\��ٯ*:>��ze>C_��	�Fu�
79�:����=����.SH˖d�ⱇ�z^j���ȫ'�A���ޭ	�V~	�� ����6u⫝̸.�rs�����R7��^Y�.)+�M�``(t(IZ>�,�F�s|���Y�2=�5]V̶��͘��8�����^��}uk:@�T��DG�B/& ���������,l6�;�};��'�BEgN�S�;`4�~���3ڒL�ڝ�κW�=�0_����Ғ�Y�/�U�"�^��voC���Ң��=�V��̞��Oz͊'-Ĕ��d�-\7]�[�����&
�arXN�h�����Łܓ�.�����0�HN������B,��d��9�����c��%f�-e�z���E�ޒm�Z#N��Ȍ%O5����3�N*�?T�#p�d��,n݂D�������E\�\��=�O,��߃��'���S�y}(�U�X�6�����#����Z�H�;�Ԟ��q�\�~�<�H}n�Xs[�"�@U��(W�	��,��K���gɕl7�i����F���k��)���q�*rdWQ�J�n7K�Z�0��x�H�X��	K�:�tv�{Y�8��:��aXx��M�&��������������D��jr��Ʈ��;����{�ŕ�X{|�U��oNm9�SqVg�0"�4�@4�G�:A0̰�;���
ۗ~z^��:Hn\7D���<E���uDyt�6�3ƚ�S����#���F�)��c�	��О0��u!���$J����t�1��?�����,�,	g��^`�X���O�1I�nTW��K���[�ײ�2d���Y����}({�m� B��S�w��Z��xS�P}Ր�1#�
���Ȼ�w ��F�Q`)�=���[��e���D$��#�����;EB�D俞ɋ�|�W7D]����"9)yy��M��������Z�@��]>¾���״�jW�j;z�K�s�_���Nr�\���c�՟7A`Js_�?ǿ�t���)�Q�\A�4[p�\�&�G V7��f��3!iZ��B���|
-D�Y���v�N,IjT�v���'g%�*�2W�'g0f����y��nxqj���]ț�取qG�	9����'ͱC�$�@����� ����z5�ZG[3��1�uӽ�q/5�BI�S��Jժ�#}m�}ቧ�����Ƹ݌w=�	ۯ�������~-��f	,P�PH��¾��L�jά��T�Y��B+kH�'�
M���"3�2�$��MI�1��h���E���` ō����0�l�o� �����V� -���5� �%QRG.荗���m���% ��ښV�uZ@_��9$�=����c���-�H�Cht��A^�p_�' �Av��u��k�1#�����Y�W�fr!yy��Ԟ�g|[x0�0�ni���~/.� �}Q4�J�1ՆF�ڃP��x���7�� $�d����.;�~''���	�tF=��%L�F��ꍑ@�J��)#cJ�������g��M��A&�'%���W;���%��_�ė�&����$�5D��+%��+D���Zʚs-,O^��g��i2�.S��- m�46@6�y[����!b]Y���`�P���8�!�%Q��s��Dq�N�\>>/N3Lh��I���nܑ�om��H@"]���"�c���:D��g͌Cq�D,Ĕ�_�X�;f���5[a+�Er�T\½V!�z�qL�Nt|���K����lHu�˶�B=���ŊK5%�bu:�
�P��H����.:��.���%)U���0�^Vİ(�p����+�C��U��`k+�\G};��?�6_/8��a����S{�^�.4�:�7���yp��˄;�(�@n)����c���m��\�|�w���:��Ȥ�u�]c?;~�<�,EO%t�j7B��{�V�?�����.!~�S�������#7aյ�m�����/ ���L�1��� ��B����e,�A��y�q�ȳ�~�i���ӣDi��wf	��mǕ1-3eP�	�WX�%و�����q���M��!��zq�@w�vs�ɯ�q�D���\�D��5�i/�f�6O�J�99�����w�?Nc���r6;ALϊ�ou�?嵓:Ƈ,]�$Mbʾ��z�;�i}�=���x��*�Sٜ0�kr����~�]a��+%�K�&n�"�d�;���ꊆ�jO��Ec�|"E���c�pZ�[;թ0*d�����LՈ������H�eK��^�I��^���<w��7u���@�a���c^H��ƚ-�Lf�&Z���n�u��O��k��E��1b�ǜf��-��'4D����F�O�7 |Шl��U|C�UQ���� ��.�?���>�g2��1���2&���O��g$3��!ߤ���%�)pY��7���G2|�w�����`�$���}xR�?3;�������fpx��O啉����|au�P|s��pNH����%��awuBm8�&vh�,p�>'���m�-Or=Va�C���%��g\E��Y=���/�z�<���8/�������t�E��@s�ͦ>�Q,f3�p��l>Z&:?ڥ��@�F���N�Q`��M|;���JN�칽�V��\?�[����Ꙙ�s������<h4�N@9�2k}j/P@�u���k&`Z����Έ�Q��ч2�5ɉ,Ę��cѫ5NTŪmy���P�'o�#�A�}V쿉f��ho7��=�;����Lzvzt�|�n�5��?2Cΐ`X����@�A��/��#B)|u$3�N�S���dC`F鑻[��dv�'������,��,��ʗ�ގ�̢��+��qQ�Ok�rk��w>�;�~�	� �~P����;_�!g�Y|;殂C9�}GL!�W�ג��U� �m�����Z�}�&	���l>v�y2�L-Yue�úk�K$�����8Cʑ'^.5"&s�P6^Ѓ�pϛ_��$�\��+�f�U掲�D�������B���'����4�33���\���]_�W�)���4�8���Y�v��2'����X�4yGE~�%�i��g7d�Z�����x_�:�2�����EK��z��u���U&��ꓝX%<�y�[�Q�ko�f�r�2�i�%£b�(����X����?�@���%�Xr�<���F+Y�/�Ŵ �UN�,�E#�Ed��R��e��N���|G�Z��k�ާ0HφX��#�W����ӎ�+)78x�=���.�Fuy$�����>y���ӂ@
^��lI|Je�.����/�6 i+G��;��ive_�S�N�\/t�e���m��ȉY�Ӆf���s`^N���>L�����Ĕ���:����v�����(�c}���?�0G�>����$^l��I�(;���%Ԣ����\]�դ<e�Q��"�I�A� 	2m��pz����_�(��y'��ke[�D1'��i��%z�u�^utN*?�ؿ9����O|�[�y�c�2#:aEc���yK2-%�HEx�9���L�p .��
�w_�������H�"X^�iفD�U�����6�6j@��1떄�J�>���� �^���T;�Z�%9��.YF�{�L�P� �u&��]����`�������lwDBaի�:��� ,UU�NݨL8��~Jn�v�ScHrTy'�_�|ϒ8y���@;O6�A$���%y�?O���F�*�qAhWR��o5mΛ��] �w��"���\���{�6����LgePϫˀ��wuh���
�rD�J�,����Ts$��|P���9�BP֌}ӳx� �NH3���%rQa�f���ם�Q.-�:�X4k�e����Gǰ���C]�u���y �AB,[T�v��Ⱦz[>T�XG˥7V(�u;�h�~9�tD��1н� ��	D�uD��Lj$� �y'����-wv�������Y�!�����-�8k��7Q0S�@�]_�!l�8�0';���7:Wu w�������N	oF� τ[X��K�K�G+�$&v1��,�]�1kц�z<��Dyf5����<��)��v7��A�&D��ܯ���Ƿ����.Һ��~^]�a��ψ�O;㛋{1����u����uǓ�N�SM�=��g���aP{��{����!�d�c,�t��f����MJ��ژ���RLt�^Z��^�0L�s��}���M����H�%�v��䗊��xc�5V>�+|:�'��B�;ikq~��Db��}\�d
�(������O}/��AA1<&��������Ś�qC����I��jy]킃���>�@^7�"�qG� �<YLt�G��g(ӳF��|:�F���l��&w�<̡&>>lt����d�!���s@VЏ�c���v��4����/=\�Y8�l8]��oB���2�~�i�	^�$���������*`*I��\w���7p
dw��&K#�J�\�N��$l�r4��:���C�LZ�ݪ*+f=ɓ�n�թ�:9id�0�����d���EH�����{|�6�D)K�K1���H�/���^e�D���	9U�\*��X4����j��҅f@�������mfj�g+%8�k{�@�*�o���n��Q::���F�#ԅ^�8�Z{��^����^�6�^	���pc�gփ<�CT�Ŕ�v���������օ�_��iҞ����/�JEWk�fma6��a��c0�3[������TnC�gh6�*>8��&;4�LR�e�	s�����r�@���Vl(D�E���Ú���W�
>۽�DĲ<=��2X��u�O�<H�#JDз�W\��l�ͦ�"���7 �C�������l���{m	�X����>ܷg�W#t��\ń��a���Ă#YZv�`��H튣)AU��ѫ�;��E�F��v����7M����t�%��Uu��,n4�A!�g/ޫn��{`�.<�U�/�������I�Ƶ��m!{gw�^��W��)����3B�R�1+�͕�~S��ސ�j���	Y}�6��;����ϟ��;�F�8~(̄��61��.3��)�H��n��$Պ�"@n8 i��|�'D���5h�"�����9Y$��!��آ�Ek!(3���/�M4���t"���2s�es�^V��&:���]�^��)���������xn/ڝ��h=D����e� �*�v8ca����%H}�r�Zuͭ]�2��b�G@�-$�t�f��%�2*��d����ǳ�5��~��o����Y���:��ǼᎩ�r2�n�7��X!/RWT7��_W� ���9����\b�5tډ;���A��79oZS�_i��H��U�X�I5�V�&�2���_bR�榴Xk}y`��=
|��V�HĤao7��/.�����H�t@ hc�����B�V1d��`�w�d4M��qg#P�
�O�����;�U�>#|lӁ���f�<��镇��K���WE��c��DG��0>R�i< PF��D����,#�x�T�x@�hQ �U�T��&]6�^7�q2Lʏ�O9n�a�����_���%�ZL���/��#&����!�~^�f�.)�����~��s�,�b˘3����w�é1�J�`���l�:��~�v�A��M���Rt�N�\A�W��Oc�pB�(M�oF��_�DeP�w�5����$`�L��ڂ���z1#�6j��^ek�~)��ͷڄ=S��r�qQ�$W�9>��ԃ��9�"�u�5�x���o���gd�+^h]&: |B�4��ܪxő�_fz�E�G����cC���h����	Q2�~s�C�H��UP�Q�C����*�Q�Hb	<xg70��ɋ�GBN��Rٺ	�sр$5S�?x���4������~V���nD��I''�H����s����j�<b�]�h�!)��d4���.aG��M2���֩���"��˦UGX�d�F�~��f�4s�}�>�io}-�b��	�ߒ>�Kal��,�n1|j�~KN[χ�>T_a�����Ւ�ݮn�H-������� �y�`{�>0�pҝ&�`�;*>?;*$C�YDP��Y���шk0×��p�$2Hd�Bk�v4�y�r�գ����Ϙ��6F24B��KJ��O�%?�f�d�P.Ps��y"c}�P�J���}w�M~����b�����:&�����5=��
� �M��h*��A����]'x�oUr�-g4U�m�m{y_�.��$62tt��Cq'<t�kb��f�tV�2ai>��\�u���o���99~Y���c���]C ���7��4E�@��3�U���@9@Mz	���Qd9*�|�.53+5�5���;�|��U	+y����W1j*�]m�#�%W{p̯`Qi����1��Ё�-)zr����p(ى���P1<�@ĸ7�R���<����s�q�Jml�&�a���j��K�e',)î�j�AS��j��Ө%�.����a��j�C؆@�s�����w�/�u`n�럡��x>�O��@��P�#��{���vy����3HI��ݘQK�C%�V���u�2�|�\����~xT�8W� 
��l F�Y�#��h.Jj�sa�q���g�H�Cu�D�=���7YU������x�j�{�S��z����6�G���"s�{7F�����K횄`�T�*�R#����xQ��z�_?�*]=��hu���x�F*�̢�!����wnYA<G�z���+���׹ѿACT��B��xhυ��������D��`K�93��j}?x����*2r5v?�`��,k"1�l�Z�L"������x�E)�܋�Ы�}� CɅ����{�q�T�H�L{S)��;��(����x�f��w�)�
��d�w�Fܶ"LY�
�t`4�M	�YN[B��+�y����݄���#N��Ri�I�*/�j�v�b50B�饇+Q���+>��of�Z3A���N�������%��flf��g����c䚊��nM�J����{�e�Uv����u�G�%���K�;K!EܙC��-�V�a[3hm=�"�LF�OֹN�dP����g�mԟiY<����E�Y��\_a����^�_� ]�{�RiB��$�Ts@+���z#$~�$,l&�1!jV��
$8͏j�{��'����u�]�o�LQ���lFJ[���+�h)�u���aY�)
T��a�?vL������� a��{jia��Ú�c{MRB���H��(�+0��k�N��<��@�\]�@Kv���W8���~�T�#���D����i�Os�	�L��M�Yn��q���ʑ��<� ��~::cB0%++�UAL����H̚���Ύ��ˮs���)�8�]��l=E�l�%�^!�g*,�g�M��Xxp���<�d�FH��H����+U�û�G��a���"ۢ�|0�=�`G���e>��*DՉ�����H#��&J��i|���1�����[�Ex�
�ˏ�|��/H�I�Y��uWZt�u����%���{�P��;�7u�͛�V�1��7�h
'u���d�4Ŷ�Ix�B��n��I�b��N�p�$O���_�c|�?ҫ�C��:8`�d��!C�h�?w�糇œ�CD�zg��&�J��L4�2n�2zXx�o��z��+�dܛ&T�Ԧ����Oh�R���9��������1�������}��/�o��7�	 �ASnV�ii.��>T�ᯝ�gH�أϾ��<֡GD3 ~}$5�)C�ߥS�N���m@�_���v�7ܚ^�d��6��J�!�93��<��GK,�鮾��d����a�Dǂ�i9�+�|hx�P����t09�ĝDZ�"?4D��M���J�����B`O]�e�_�].��d�+H� 
�:�4 �4==�$�
�2Fcq��}��vĶ�P����� �q�Ǵ�mO+������ܳ��oV���Ī|7qT'��휭ҊM���v�Ѳ?��ug��*jh��+����s���ܞb �C���!=�U?+t�ʄ���6H���?��?$)��X�B�'4��ß�����^-g���`|��X	[V�~�Υ})k.�-�7��oL�}�\끾�cJ���c]x�Ә��9jw��ԯ@�uDS�]��L��G}��s<��F�����֡o��)OQܴ���@��8r,.���[M_�M�O�Q@��mC��AHhHd���S~�&�y<���Ͳy�����m�D�$"����Y�f�R�GlJ��z'߃���Y! ��~WR�х�GF%G��F筣.�֜KAѤ˔Lܡ�p&@U��_��&Ƨs4d����4��-=��Pal�#vLޗ�ْ(Rlw��y[pm#.,�4�qw��E��9V�E��d�2��2=�K ��/��1�G:C/���q
,�cqI�$u��
mZ�LY��yi�F���~)���>�Qy���������6@��W#���<�{9m/V��p��O��T���/�2w{�AL��0�m.4e��ʩ(t��`Z�	�!��$�ݻ|��%1纇;)D8}A@�'���Ap>+�.����>�{���]{8P�*�����s�� �HԈ�kO��Õ���Q�>hO%s��K*Nz��Ր�ӑ�΄HU��V������=�K;��w���d�'�r#�T�����c�T���<�z8���d�h͉�����I�e��L�i�a��;�#"X֯�Gׇ�N�kӭ��n�r�"K�m\Ԓ�L�nՋp,<s�5 ���x�|�j��%��4Ɨ�b|�G��!�@�F$�t��[g�飿2��a��:iHo!����$q��a� ��y��8��v`<��|�ybt$��J�NH���kL[���,@),ceu��Ƴ�N:^fp�?�\}cbX�2��J�f$v�s#}u��#��_|7oq&��Rx-K�Q�����0���uA���ͻH���cǕ�Ϲ^z��!r�-���NO��E����\������)��j�,���Hת4�>�����2�DM��C��5+��2)������(����	�1|zї�e��+Hy^��B`/��tt�-^�M���x	�?�
�����'(��� �tt����B�q����5a^!�_Z(��E#�{'�%I*3�0����H�����4�������l"/<��kK��Gg��D�P�mf����@�I0��I�_�S̤r��V~��%�����+�zh�E��pZ���"���۽��p$<�K(�Nu&o��Jt���������n�v����KU�~���?c�`�׺�/2e��� ��͖�/ i�_�AZ���x�z?TI��"�<�K3'3��87dè6���v� ���e���2ϰ�m&�&F�C�	��,�뻨RN���1�a����}xB��!���}�:��I'���瘒��cCƍe�����_�G�uyϰt�E�VA��/ƿ)W��g��òG��ZȌ;��<�'d�X?�ζ�Y�ܼ�d4�'[*���iy�u�@�\\��7�����I��ե��2�Zv�j�{<3�:��9O���I�����֯�sV�#S��)��$�-�n��v��1��V���k�<M Ŵ$�#��2JizԎ8�1)���c�������M����������&̰��I�Z�n0��uS�33�ְ�A� %c��b�@ݨ�I�cC>yL&�09E�;>ӊ�&����ѭ�G�Z���c%��X�a�ZFr-��c5�%�l�t��4�e�,G��lF�;�Ȫ��]��^��),�it�in 6��$��{�x����ìsǕg��Vgd�V��_و_��7��Up��9���4l�W�a�b�!�O��3���@��D��)l����۔_�1�A�s̀����7%�fꎑȪ��:�[���M�\{�&J4���yh�����B0��cEK(�Գb��/��`<�~>�7逴�ThJ���`�Z/'�$��⪑L���sL\�3~i�� ��b��j�����m��عe�>xnw@Ѥ�c���'nS�w��%�}��a6k�|� �yk��x��e>ٖN?zQ��*(�pX�'1Eʹ�����n'��}y:�!��?��G�/z|ؗ��E"@�s����>�s	L��Pl����n�4�$�Zo҅Nt��.BY�8���%���ɺ�0�O�n%n���jz��`�9O �\س��|��]��,�9!"���v���)+�����l��eh���	�Z}<@xL�5 ��\��y��9c᭚�O&��k�J"�3�۔�O��{x����xU��T��b� F�.*:^L�m+�M�ֶ濕ږ�`��������]�/ ���,����ҟ�w��q<Լ=�u��ܹ�ݷ�����)�s'GÀ�E�G�o�~�u�WT+Y�RJ�Y�B��D����F�g��r�s�)� 75����ϬY�̼܋@�;�#��t����ĳ!��ҺeF�/��uԵ=C���򲰛�9�f��t���]g?��G�v�����tw3<�����s��TB���{�P���U1�e���=�:ڄ�G���3�&�쉊��3�h�p2hS/=�xK�o���<���;�=�ʕ"����-�c8<���Ӻ�,Tp������?�|o���^E�����1����(	*q�ЫsD$��[��x���%?B�jRqk�Sh�h(��g"f҅LC�])I����e<�SSMZ&+,Z�{>�ڻM�(�Z5�f���aO��.�/97�������b:�?H��5Z̴�@A��C� 13�f����F����aP4�����(O���i�%t>��&ꪗ�#��1X�e�WW�ʈ����zT����A��	�ҏ���&������,�镡n�o+T�%��T�!*y�"�(YzX���:g<gCޏ�o�;\C�Ґ����]S����H������!�VN'�cE����� LOh����.�ڤ�{i��e�E�}8��;X�V��Vp� �9 6�:�0Ѽ�	*[�����a�AG�\�ƀ55'���	�8�p���kA�����,{W3-�]|��jV.���K;�#c�a6�Ή 8�j�,�↷	�fnY�$tˇ�/����k&��Č���"�m�D�C��*bͯM���*म�ؚw��-������T��0��&�5�"԰BK�0�L����e���r��hg��p�b��+얍G9�;�V��q�և`B�e��Ʈ��YOǝ��o�s˴��"*6�R�S`B��E�g=H<��;[WR:6qJ+�t��vY��5z�:��5hP��f�8��1���;|A0	5Qk�"���Xn��c���W\L67��H�:��i���5���@j�Ԓ[������a6,* `y��L�r��T7��Sa��ԗ����B��_���1߇v��=�LY\k�U��]�K�3#+��D�c�����D���x��-�[j@���'�.�;囟L���.Uֆ��*6K�ͧ9,h��[N�׭ro���՜%��&���;�@��9��J���P�G#����|!� s��e�ּ.�����R#�Fh*W�Xx	�N�	�|��ɱ���<����N��*^/,V�~�]���Q|m[rl��Ў~�/�4_;Koe��e�2d\�!z�����DF:Rk0��ɳz��=����{�4`���#6����57���z0�W�]�-����k�QK�9o�tn��^��ꐵD���2�c�zL.��;Lu/F۷5�C���H���5���ե�F����Re��ϗR'���"䲼4�-������xC���S!5��-���M��/� �f�M�1�}E�BHc~��Q�tw�(��y�lWmo����Pq�ܪ%����iC���U8��y�--P���	]2��N���oq�9�̹����&3�_�F��Q�c ��{eh�Z~i2y9d4c\#��
�E,׭چvp\���h���A�B@n�E;�����+��1�8'5�L߽PM��zX�r5|y�(�Z��ec�:hEl�^4����N`�ai����Q����ph���R��`R�̏p�܌z�֨@���KԒf� AZ33����:e��*#n��/��Փ���<l����8�߶W����gz�'�<��.F!��[$J�iy:�Kg�@���{�j��0�8$�#��(e�u��aƢ�M쐳R��D�y9 �O�.�ȇ����Sn6�2� ���6>�����3�;q�Qtl]2�'�s��D��E�`y�V%	39��QƗJ���m��
u�܎F�*0�9$1fR�^6�_?L����IFoq�oj��ʏ6����$Q�{�����<(����R���?=�^��!��D��B������J��i����q�iC��x`1�v��b#�L� $���mw�#����/+�ჲ�GN�����$�V���0l��^&B������X��%����h�+͗��y���N����D;���v&�a�n�FXA�T[� b<�o��	�|E�y�97'n艘�.-�Ϡ��9�h�8��}�E �IP�0Ɖ��4F�X_q���+)ހ�`5*��*��=$	�^�K���l�&δ��[eI��p ��Ha��a��J(�*�T:l��˖�
�۶B����Hd@��#	4�{.����R��ˎ 4������6fd���{�!د�L��b����;��C���-N߰�#�����`��yRXk[W#IWWX�%"F������Q$���)0��*�N��3~HȺ��*拂ɶ�~�fn�e9GA0�z6�lvS�Sf��%��f��g�>m�Bc^���_`�� "ǻ�o�(v�m�~]�ݸ�2n�J��O�[�+���e��X��R��k��#�5n��9q�d���JѪ���X?��V��5��7�ū@t�3X�;"��}�z�ZхM��*,?����՘�X�N 2(�%���L
������fyզ�{e�[��/��?w���/l,�d�0e���)�QN�|Z�b��6?_4�S�V���@�M�ɉVܥ��-}� �wg��g��Ve���Bb�o	��JBݺ�8K?(�@@��Q&��o.��%�諛5��o���c��V�ȓrge̷�h��-J�ѴD�ęJ�����b!�F�$a=B��j?g���S;�:�ካ����ld�r��1�CW"��׷%�9{U l y�V3�~��a�����E�$ܘ��y����Lqk1	����P^�w�2�)�۠�Y2���
A�������I7�W�8�$�Q�~ub^�/��ɯ�����e�d�8}�8��R�p�x*&��{@vZI![�z�d]���vش�O����)��vٰ�p��E!��y km�P�+��K��qW�;ط�c��00nhյ�P$V���4�JN�J���e��D�7f O{��`C�L�7K �;.&j�V� ��t�����OΝ�+�d{@��@s!�6���t��/�l�ذ oYig��>�K2��-mJ�������zШ�b���r��roz�橴)D�f��k�j�z76�I�d"�I�z�o`��#/���>`��y)���-=%�[RO?by�:e ����N	�J6����'ubE���Lv�l�:�/G��6��<揿����:�)�0��1��Rܯ*�t�#h�
a�J�)#oJ�L��BTu�/x����4p ���i�/��3�׈mua:��)u�js���g�v��)��s`s�Y^�wb�J&f(ne�V����ϭ֟���� ��wæӐ�h~&�_��w��J����k��G���e6 �쌉�9��'�p���D,�	�H�\\�8=����Rk�E9L���$l�����g�u>�3�'��l9�! I[�}��k� �o���@V,�g��1w�[��!�Wƫ6�1�%�Vo�y��������?��M6�E�`��A8���W�fJ���4��0\���่yb,5c�ѴW&Z�72j}�$��i��$$�0�50��������\"��5������<ҡjB��:��d�kE��k�J�h�}:g��V���FL�yT�}���� GD!��(�;d��vC4#�?��'�!���g���*ڈ@�f���������Emu��5;
����r��.D�,��:N5���ʤ�1�v�(��?9��cP�.n��$���AJ�yV��^���#��~��G�$p�����G���п���J�_W�y������^*�������pYu���pf��.�ω=�ueېM)7�F��gƣӷ��sYd��ܽ�}�{n�0� :�F��2+��d>�1dp>���ߵPtr��T�Cd-�J�m�D�4#=F-��0N2@�
�R1
�N��R������d@Vn�����a��*���\�I��)�	���G��M�(F�����!�h���2�_��$��'��c�?%oF�����C�t�`/�ƋE����ZxG���D!w1�Kg�NGk���6~w`�(�9�@�Q���<_C����]=����%���ǈ�<�R	�#�\�5mJa��dbW��>�l��)KO��t�1���acc�}�p�K�ɮ�IOP�@+}}���<��g�Ե�3�_&���?��;p�^z ��lܔ��\e�S:��%R,b���#!��Z��~��a��ˌ]Y��T��Ns��f����cXw������' ��6u�*���8���6]|��.�L;� i(hX�1܆�����6|�y�6�$� (P7u����Ȃ6߅/�^ޠ?GbWi�͓���J-��d�I�q¹e����6}�:XEI�G�����t���~��������͚�ӯZm����؀#�ȼ.L�HS�¯9�T��*��8Y+k%��٤��!���N*�Is��G��et���d���Y�F���;��vdJh\��ȑ��hQ#�<�啟̳�'��bD`�i����:�?B�⹁�FѝDC�\(��>b����ѫ�B�
h���b�trSyE��^�ҧ��>$~�W����D��T�T'�^>wx>���|I�J�j޲�H�PЕ��~��ڗE_��pl�8:g�.��{uX(�?�bB��gBD��!
b��Vv\ȔG`/�N�2���ru�khnj�IǋN��#9fy��R�H	���v}W񪤏^L��ƽ�ٛ���W��&9�>9�U�$�G�nhM%�CL�&o���[�Ũe~�̷ �c�]q��#���P(U������M3sV�{p?f��|�HM�������I�P6JZ�t��U�� �
~���M�^�yPb�X�)oD^�-:{�9��2��k>2��"'��by=8.{�h0���� �L�,����g�<���"�Q�;�ϴwG`��X�Ŀ�W�����$A�qs;ϼ��p'3)\�E�6(�)����H
đ�kE޻�Ig&i�����0U����<�U%,'��c) ևAC��(�3\a�S���2�7i������=�"|'�R��������Q��nA+��J� (�f�ø7��b����@z��Y$!1z��5<�z?�I��݁����m����,��A���F�4�s��cL���g8��xP���NQb�9p[�K�G� P�("���[��l���
N��d99�91�%���p?,��C��Q�l�\���U��,T��m��yhgt��_��;w��L��]�E+�ׇ�+�>�4s^�M3�7ͨE��J�׍RW2�߁B"|�	k>�������oAu���x_��4X�0"�x)��-�}�b�O�VU�T�tV����+?U���G�C�.��I�y�3#R�c�npy��OUB�tAE���/M�A�s��3֢�y������]vLnJ�kE-��	j����I1�ђ�?�:���k�8K�\GLa���i�E�6�G�/:�H��#� 2 MSa�>��Kp�؏�>Ӳ���d�fXf�L�׉���'y��߆]�T<:
��Պ� ^��p����`�m���h}+�Q�Z�6T/�qƏ���)��o;��S�܉�.���f�U����D�pe0?x\�e���QeE"N
-�O�����鰬���Wy�V`N�s��j�H*H�<1����`T(�JC|1�{b�AT��n'"��{� o��G��j����h���?_?��rA��}�m�3�W� S5������4x	7հ��q�H�=��(��b٧�<����?	G{*o�o�$�%�_���j�*����v�+/N�B�;E�@��C17+_(A�[2�iͫ��:���H��D��{�w��~t��_��z�;p4�W��8�k��D�? =Î�F��_��?�v���0y��1�.�l���*�^.�xR�a�A-���9o������TY��(�-���I_m��}�����0�rM�6��v�";�y�j.�r�ƣc���x!C��v.������~4�w=���_B"
�׵���a�3���M<����lqA���w���C�ίVl��	�v���F1��7�f��'�b�߳��lG0���)�j*τy�x����Z<���,ہ��] �	�����b���5�?�~��vX���]�o�%>yc�H�Geʌ�	^����?�q��m��)�����>���"lkQ�]9����dh��Ć9v��~��]����S~3�7� ��
�j(�b�Z6'�D���a��Ω�#yNr)�����]O��ir��	�}L��� ���DB��`��Ô�iC7���Tދf�����TҜK�qOԚ�>.�����P�5�vD*�H���sA0�"�����>#e*Yn�J1�y����/���qq2J����qR\*��<$jg�Cm�iJ>��9J���E-=-���(9c��CT�gO"�Ԟu��ǢTB��S�o�E���R0!��w4�)%�"a�*�����?��~��e
�x�<��x���AN���_��AK+h��E]n-Q&~{}�o�� g�ZQw�v/ez��0�n�Fi�JK����קoFږ1�����kd��=:@�W� �����;ϼ�܏US�و��`;Y��H	:t[�~>�����S���9����vH.�8�<.��vnH�{�'���8ň;3BAfMj?FoH�C�Vy��#,#헐���a�X�h+U_��d<$&���MQkK�$?�R������-t8p����ᆽ����cG�e|�4^����'�Z��ǋ�]��7'�q�|�E�>_Rc�{�����¦��FQ�t��Wv�����3���L���j�?B@�!�Ε�O�Ӓ�|�R��x�ԏ2��
����[�ƴ�<��9���F(��exR
G���@��.�������l@&���K�ulQO�`_-m���7�P��fi�zՇ�5�W���gw׿�0r��ф����������RW���e�y�R�@��)	g񭑍�:��U�L9�b�7y[g,]5��P�K�k��>�h���jԌ�Rv���0�o��W�4Ҳ�Q���	��.k>�Z�G�ў"y�9�������0��c�vv�hiXn�N�_�dF�6v����F���g�oG��뾒����`�w�M���ϰ�'�;�F��l'V��A�9����ͪ �%���f%k��fE
�`+]��Y�換Ș��gp}�4$kq�ٛ_X�!z�O�0���G«ֻ����T��Y���������U �'�ڌ	V���U��di�yg;Kйڬ�:&�d8���/1
-��z(�y��� ��"O�*��������|�J �M��@��ƹyjt�ved��l�k֠Á��.V:�Jw�`nX�v�K�~DF��4�@��|�x"
�Dv8f�[�|��L.Rz�_�wϜ��Y:Dbd������9d���`�yTޔ�պ�q���v�B�(��,p��浠k��@����\o���k��	*.�np���MA�b�c�)C��/Y
߯q���u�?�C�����8M���OHa�9��v�'�hR�^C]��0�[~kSY7�q�C��(�G�=Л�V��;T阭Y��M?����:�%�j!���&y�����1������i�^�,^c��qw<Y�H���%����h�I���M1��H#"�e3I�ʅ~���U�x7䤤��\Ӊ�����^�ʹ�p�Q��o�z(�]� =r�Q�=G&���[`Qy�(6oZ�(��/p"�nG���I6�Q�PB9�_$H�l�S��?%5=�XY��N.�&�Z�L#8H8.�.�t�f�jL�����_I]��[�L#�^j��/��V@�6�-�����MVʍ%�tr<bm4�G>2�`PS�ݢ����	t�4�x����� ���ĳ��I2�5�R�%����ps�A�B�(�j[�NӴ2W6�?�
�}��` 3:�����!���D<S��ߔ����w+l	��e��ᓈ��޾d3iD�!�wl)i7����C�lkV�Qvbۺ���5@��i5q;nrM����'|��Ԯ��aV�oD(��"Y����i��5�^F�F1�ao ����%殐�]�9�qz#!�(>�Ë�Y�J�X^�� �V�F��ž����ɲ����������둓�B���v{�
<��,ѫ5Ӧ�ސ����3�g.� ,��M�x��R�G�d�n�;OD_��C���.Y�~u�#��rAo`El�b"06#��(Py�*�RUjdSS3�k�w��30,� Aa��������Sg��r��)��}�?㋶�O4w	���Tb��	�+v�W-��^2f �G�L|>�wy�W���,��=�Cr�Ҏv{��i�6=��1`29s�_$� ��;�� �)�T�]��8^+���NNR`\O2���a4�		s ��ld���4�V����@�����4�іWO���:��F���J��	m�$�-��b羒NC�ċ��H�A�w0/GN;%�U��SxP�7P��G8&`Z��_����S�&�/o��(:���-^s��+�.���YvY�k\���]�����H�R
V�v�:VH����@b�s�T3��1j̷.e��د��� i�)�x�0�������}�K7Z�j���>��U��f4n��?�V(�P�r�Q��G�e�[�&�B��In���"��K��e��:dm|� v%�t9�v�S�x6�̀LUh0����F�~R��.��ep��e<6j�,�/J�ѝrÑ�o�/�D!���4��5>:K��xd�$���i
���8a�/�;�T������ӱ��q��~S�uԫ(��QyE��dQ����jЀ	.AL6�Y&�~�)/ݫY���hS�=Ig��@x��) ]G}�2G{�J�|<�iN+�3��ߝ�Nכ��~|�_��X��X{mG�{V��Jk�p�s��~/���θ�������B�ۃ|w9��|g�U��h��꠹j��}�_|�y�̏"J��fΡ�z��ք�����߄6:� ��=7h�BA�����r���Y08�$�}B��:��97
�[���ތ�dըѮz�Y���D$뒩;u�[Z��Sݴ�]p���%~��oQ�ޗ�d�8Ŧ0M_Ƿ�ء��ʉ��)a�8�eK_E��&|;V��H��,ڕ�y��<�z�p,K2ض#<8���08������*}� �*�`�C������^�q�qx�$]��
"��Pn�Z!�eA�l��±n�7�������vb�v��K%\�6BıĔf�6��/�s֝�d�-��/1<|$}��6�u^hP�����O��M9��3�(f��ևb2�H�b˜�G7XX�9��W�ܓ�R
3[T�Z�@2�=�eQ�����I��������;��s�)�������dc��i���Yѻ%k�P�d�]�H0�]���<P?޷r�u�ed��_^{Ny��F���"(誕SĴY���4�߲:x�;����;�H[������x�;�a��D?����c�>=;#�tk�U:d����Ќ���{����9l��܏�aS��9��N�����A�/�X�>|�(�yD:�v�;��R�j,(�5t��u������ku�ÂκS��I�~�K�Tp�s���r���JE$忓���"<��?�*�}ZM�v����w0�n���GP��n-����B
�d���M��7΀Y	 Nڛ����3�.s�!{�k]�ć�<Y��5̏c6�|'�#��~�5���?J#�����䅲�CM v����C|?1٤���;��4��b�6�A$��%U�rη�}eN�u�1��>-�k/rr�U�3�[�t�� �$�_�nd����`(D�5�怆)���А.E\�S��^�!HK�L�-��eY�Y�KU��fJ-���0�@$9ޤ�Ix���z�4�U�d��j��0�[�����0g(hj"û�9�W)�{�5aE{�EPg�Ę%2�n�h��2��g�I:�A�f�d��C7iT~Z�	T�o.ۭj	<8-�Xi"۠�N�1��p�	���
�%D�&�~�ο����:�+�cdZc��k�V-��#p��%���n��'wr�5|h�F�� D���)�V�����j��[�r�=�� ��n�(1ԣ�0�Θf�L	��w�V�C$������t��P�� '֖��V��[X�Uɏt�ǐ�_���d��Aᬝ2H����~ۦ��`¥E]�|��v[2���B��K��I�H*�UphRP��a ��e��l\���UQَǟM��)�E��H��/�X!5�.{Yc@�㐎�+��txK9�#/�,lxPƗ4,Dsjc}����m$%v���oC��
	ꅣ)��)�d�c�t��5�o�k��K�rH�O�c�2br�8L������S�Q+���wZJ��$)P��M�/$�闽92yC�u^klZ5��K^��5��@�>W�gt�4=v�A@��Y��P���)��B��e�[��U�n�)Х�\:�UUt�n��E�~�O
��e~O��C��P�=��������9ߜ�`�-�[��tQ��aғ�CՎ�G$|�\�3z�a�^e�\?�����+��@�
��ۋ˥~C�/�nV*�\�����6Q�¹|����/#�p������*UZ�I�d�־�0���N,S��J�m1�o��͚�p��,nB���f7���.���sx��󙜴��� H�!�7�i@��z�aP|�cm_�	���e/������׾��4F2��Tw�uB��f5�TG"�.����X��<M���c�/��LdW��bVj�}&���b�7�~V�ۢ�m�T�֐]����(�<Vؐ)R�֠�A �h����4vMT�F�Ү��m_&u�����LGiZ��>1�a �r�_��^7=ўZ#�c�ސ�����Ls.XO+_2A!Fq��%y�����L�S"��tu�'��k�;f]2��64�
��2OR_x��#��|N�օ���Z8[��>酦��:�cC�V������Aq?�����ȷ��q;��J@���J.���� �|��<�}'d��-�1q���E TAk��ss���H[��C� ?���fv�1W���<8��g�:�:T�]o�if3eD���)g��s�{9IR��[|�c*(�xp_����qd��Ӑy�3IY��XMר��!�Tz�%�g��N���A����Q�t�r#L���T�:�A6&utP$�����p��54+�X�(ZGq���z��~�	Mc��j�\C�B�4����VT�d��ޭl�u �ũͫ��>ј�}������4�}-�����S�3��K��sm+���}�˦O�(D+W�Q������鏈�ٴ!�yZuFA�AQ��)谣���ڪ&��i�D��$2U�ynQ�1��`ƇX1J�+�'gtV�#8�Z$�$缾���8Q,�PyF�S�ʗ{�%ۊQ.�E�y��j��pW�*�ٖ'p``�.��>tctf�b.+8��A������cX�WT1�Omٝ���E��/�gr�!���%�>��x�~��c�̽�;�7���v��������(O��uIP���E���ϟk)�d�m�KE��f�b�-��+�����QKol�'WO�b�[	O��y>��X:�Dg�8L�P9�\��D������3!�%,\8ػ\��MeGbZ�G��FR��C�e�![�V��2��I���K�
���1:��` �M�86�9̞� �W�x�L��w�Bw�C�
��$�\G~�?~#*��y8�\�!��w>���ǘ���x@=�*D�����/׫݌�}���8���y��f}z����F* �8/q���<���O�w,vo���c��+�f8�ǈVO/sH5��Q�Ai���|X��
I9���G��2�穡�8�%������gCŶ6G�db�Od��x�2-�Q�缾x�R1����E����zNQ��f\2�S���re@�X�����I|j�H�(�q4n?���Hp�10���� �Z�n0�e��u�齰����rstp��ƢN�x:{zB5�_-���-�����F�'nY
���:Lr(�24,�8|6VW��j�ˎ��7����˺=y�*�Z��'%�$��{�eșXsp�9��Q �U�b����v�pS0ɯKp�0L� ��L��:���?@�4�3�p���B���v�$&d��l���}�>(��;ڿ����3ŀrF������_��J�رE�13�^�¿ev�vd��~a�Ӄ��=f���P�+�[��̛E�(�rs���Nͱg$i�.��'��r�͇y� "1O.�8��}�"���X�k~p_���-�f��ό�"�!�!��pS�����G����J��!�l������S�������Cr����:DyBUd�mp��<��b8�DdtI�c3tu��ܺ0������a�ιX���b��׊�9�.�7?X�Q�.����/�����M�3W�Q$�D���<x����Wcl�܂�r���J�����U,1ɭ����z�$�m|
��P�ʜ��A7��$�����?�nޓʍ#\Vr<m\�l�G�.\�|b,��봏�.��w����Z��Kc���+�JR��'���L�E�[��_�˂p��i��K�ɐ��Y�H0ݘ�m��6���!��!��O��)M��ɱk9�޴�K��s#��k�5)�[����^�渠-�Pz���O��;-q���]�_�� �^�AV:�LD�yN�1w��M)H�t!=��������d����u2���IZ�O�n�U�����,�[2Ӗ�!"�#)1C�k?�11�hü�`��\��ΒLI=����"�H�-@�ܥ߫u}[��O���G5@[�PEW��������!W�@�h��Ǳ�eMD ��'�����c'pxxb�\�������<B�U�Qf��E�^o��]/���9 ���H��4���6@$ՎT߻���l��ᶎrZ�K�*|s5��>�UT�����'1A[P��§�wᠣ֖�4]`E��X���t�&���[&�y���*�:V6�=�����&�N�ԝ-B�Q��RAL܋O�롵�+&S�O�M�a���\ٚ@�N�?���-J�K��R�P" Ղ��R6G�sF�?9�q��%�{�a�<�"���Ü�z�Շ�(�2��BC���_s��&p�q�7,�E�s�/�O��6���pIQf�o �>$�D��i���G5H5"��½O��w�� �3QS�ݙ+��n![N��T�\�L�jh�ݎ�<��j7���s'z�As\�>w��"���I�m�v�v@](]�p)��"���u�oGY����(��u�, ���څO�x���"����GS�B83��}�H��|��a��ή]dM��-��S+N��� *5��a��}�Oᘤb�?���栮~�����>��Wr�ƶ+jd7��,�->P�8�����kf�!fȸ}��j	w�ў�'� ���|�B��bRf������.�ʽ��\bO3�vڜZr�;�c�5h3�P������dCM�5���Sh�/�D�������&�bR/xf4�M���i0�
���|�A��q�bX���E���EۊYqa
�9~D��:�T˾v<�`��� j �O�R�؆=��KI�7yݬ�AL��;Ŀ,�._��rD��NS�-(>��ڶobxχ�y��]V~�B��})��d����n��nOx�Ȕ���m\�aVj!h�'|b"e	�x':Xpo�).���%[�Di_�*�@�75K��Ļ~��C(P������l���~S�s�˧yT{3���t����z�R��utI��Z����L�x6`�;δ\Q�߼a�74���9H~��]��P�6���,��$jʓ&�nti�wPyw�r�X�~s	#�qs��7��H���w�LT ć�^^H< č�)�sG�+�V�^+b�I/��ŉ�Vɩvm��{�IhB�k���!��/(}�E/��D�Eu���7�� �x��
0w[n�Z5��̀y�7ϔ<G7{@�ɮ�.,I�_��������V��M�{Г�g<�9��W�s�� ��:���� �Q(�us6i��H�fc�gJ���W��ض�hMe��9_�E-�� �/���V�|@>?�N�}�ҿ}�������}æ�p��e�=�1I6���jO�^��+�7�p��f�}���LUwǢ	푁t�l�AKQ(�BW'�hd�cg`���r�NQ��I�#	��,O�op���?�I�	�l�Ոhm
�-��;k������r[��L��W��Đp奸ʖ�r���Q��mrB�*�\q�q�1[Ԡ��B|�p2�e�� ��)�B�N9�q��ˏ��߽�,����v�5��E�f-������wF����%�������W��w�t�,B�N��ؾ�s	O�o��|$�����i�ނ|��{m�a�����N�ؔg��hj"����U��OH�|�v)O����F��!	ڏd+U����<��Rw-]Al�@�'�_vM�x�5�cϙ����<ȒC9z0���Ir���!�ŝ�k�*�ePC`؎��*�Q�g7_?A�;����}��46��p6�Eq�52JysGp2�k�w�mF��Y$��@��%�[s�َ�%�3cUR[D0�4�Q�t�֪oP�3�_:�ͺ!�C����F�>EK�.��\�*��s:lg���:��a%�,/h��Y�;Ue6S�~B0~��0��&��\r/�0��^�y����xJ�䩩���P@{V�R�]B܎E��Q������U�3��ݠ����b+}`�����$�n'��'3�+S�~8c����.��(�2��&>�f��L@n
�g��v��0H��lZ`�ç� (t�d��Y�\���j�0ew����0
	A璃�^V���-I�����	��/�5� �Д��a���(���4� eQ�o((�{��q��U�XB�sdՍ�\k��^�`�MD㊜Կ���2�h���i[�gk�'�U،�镅9�Zvk��p��W����>F� BL/@c�F��%��E��}��o�R�X&8o#���+2���6x�n��:��&{:|SȽ�o^�攰�;jG��!���� ��ot����K����L@㾞���}8F�
	J�Ķ�'P��
�`yN�˔B�/b�*	�&1)JX�k�u�/Zg=�8Y���L���c�x���I�w�:[I��މqV$_J��G�k����#����z�` ݺ������%;&Y'��ߦ�l�c-qj��w��on V�Ucp�x�����-+~�+W<tBFEG�
 jH��8G�=e�~n�0rVT��- 3�$������{#��d~ߌ ���ϔN�`�Wgc?�:��\
yHy��U�z���p,x���R�IŐ߅J��9�#��@H��w0Ё7N�"f�n���]�'��x���qR�^�C�Y�����9u�׆ ����!=XF�,a�n�|PB��~��!��-�7�አ���Y��%��z?�J{o�m��y�Ù��p ���/�;�eKN�X��rA)Oq'nq�2B���������(�f���d	I�=4��;����$�C�q@�[��ݚ܇��r��������{1�'�9�g�T���+�4�@�� 1�
���FM�>L�!�z�����y�bHuvB��&�.�"P�N2dr8�r��?���i���]%Z�XL)�umE��+�,��5�W�n"�܏}�Bc�̤�
Ͷ���ξ��HC	Dhm=}�'���T�j�)Y������`���i�U�F�
u�5��=�]*{�UT;_�Ʋ�̆R����(Տ�^� [�D��FV`�����\1�|��'�#�q�Ph��*u)'Q�̃�������;���?�w1�"�QZT��Zs�2��DD��i����-7�Ȳ��� �PЧ((��!�0��/�u�������8;`E�G֍h��~p��X>T��f�Z\�{Snag�v��0 �`��+�%��!�j�Ԃe�6
-XŸ�($��5��r�oڙ���0�����B*i�� �/֮����"~Y�r�CY7�7�P�lK����5
�,���b%�������~^;����.�/�O��4�ʝˈ���M��Ƀ�Wf�Q��m�P2�� 	]	�����d����IM�N����a5*g4��-ML������3q~͆(��|��4�ʿx(M���0!�{p�ܚ�3_e��
֎��-�ﺖɮ�&o)�F��3~�9.�O�m�[.�o~z�m�3-��S�Z����ry^�i.�x�<t&�g-�J4���x�[͝��`0� r{�t�%>;F��X}��q\�[����	8�����0�6���P�P	�w��u�E��/��wp�u�hT��DHFGl(�����5��.f��NX~�r�U�˭���M��+)C�������,�J�US�Ob�FL�隢��A��MK��k�_�U����t�9�Uuv��G��e#zC�
�b�?�R�{%b�!�lˀm�&.3��N��N����[b꿵����I� �%����Y�$�1��X*�Y�7K��»ʌ����JU,�$]֊�ѡ�<�J 5
�!�^o����)���qB�Oa�P��S$�
�ǐ�}���%�d9��ލ�z��ْ���Rb�Ğ�E�y�l�z;�P�?�0����C�b� >eK"΋���ǡ��R�k�2�Q"�.����AT�H�'�����X��	)�����0��]A�)��m�[#�X+�nuV���=|�Win"(�趃����В8�Ot�F{���պ�[U�~�%�%*�Q26��?")F�S�W������qE=XE�^�{�~�}��@��~ 7���R� a�	�^%��^wOZcG�o��,P�=n�j6�#�{P
=��ƞc��S��b+4�ޏ���:u�X��rQT�[w��$�IY�]�7ku�"TVH�Sk�Ġ6�''��B�DY�������&�z)��V&�0M`������n���%��k|��v+�
/ϭ�	��k|�z�t/��yG��Z`��3SN�dHЕ��>E�+� �e´��9������i���f  Z@z���x��@�S�fǉ��[�W�+㥃ݘ�B99#�k��P��Q�"@M�R�(�=��m�˗��ы2O3�^/�j���g�b���ۭ��i�7��aWx� x�p�,���	8��.\�%A�{�o@x\]��"�H�T��ʋE��	���s�?�14��X��O@?��D�g�B�M:�}�߯�j'	q�Os�S$3�5�}$�&-`�|P>j9�|d�╝�a��%��!o�<��oO�k�_����^���y�0�!��͘|�۲@������;7/��qfgB���e��u/��ĳ@NC��������b�����h�2���H��
�H�C@��x��2�oj\2��(��!'ĭn|��|�3I?�H�}�Y�������6�x$�uʠ�3��$�S�	�_D3� yt!��Ļ���,���̊���W�����,j�7��Ӿ�o ����{>�3.���* ��ԄM�'����I��b ������^�?����栛&n���l��f6�A�ȉ_�8��Wa��v����PBi��=�T���26!����?̪T��2�j絸z��"�	`�H��+��-XJ���୥��(�wu8��Ew������=Cۢ���`S�+�o$)�1l1o'H�����o�������|��ܱ�D�ky���e������S2ccK<�]�pjiϵ2fO�C�Ȣ��Q� ���rmSz莀>R�@!.J����q9�PP�L���S}E{��v�4�U�0$+tS=����ճ~ⵕ���w������!XPe@�H��v�98�å���_	}�g���:1�~=dJ @����,�_^v�
c�Q�s,�!m@�Vi�N̰��E�@�&��r������0�d��2��FL1�Fk�ξG�j|"�]�V������w��\Ky�z���,Pw���q��!�2���3���:CȳP�S��5�CGL|��lL�s�k����L~�hc��W0d�7�
��	���)���m�;��V����!B\U�0�i��A����Ad^�6m�B�Չ�Ν�9���_~m8\�@���h��%����b���X�#��%7�7����	a��E�4}yf$G�ؚ�sB}�\�bݜwlS���N���M�jZl�YGABo&Z�;�w�8Oa#f,aR3��V��{ڍ}*�;���A�-�f���\��e�u@o�՜g"�����o����8�Q��:�K��H]��c͎�6�w�)���F�?�b���l�%������sڃ�-$�*���3��n���'�Es)�"4�z�d`W�Z�ÕC5�@�q���(��;���͊/$��2���þ�X��I��ޠ&����p�<���Q�a��k�9�#���o�bTnq%(Es��u�(_>Ũ�&������B6����e��]�(y	c�>bS�'�$L_��"R�du�N� �o���k��XDg�Z���θ�6Ӛ��SN�y���G�K"˥��sY���J?�nM]��<�.j쯦�چ�a�\��e�';/{S�G��3��K�H֛,�9-�g�N�v�E�_��^ҋP�]�g�Dʎ�'٭zO�9�Cf�U��s��
��Vv�����W��� �pi>\�QX�/i!.���K��n/���_�? J��ޭ7$�����O��`�2)��9,�%'��iT��].�m�R�t[����dγ"�ш�d"V��%�
�J�k��hL����ܘG�m��p�TE���0e���Ug~�p�����+��\��Z2��$x�2���[(t��uS��Db�*���Uꥺ�>#0;�O��)F$���8�r��E�<��Vg��L�Sh�N�����P1��՚ri�֓G�`��tΑ�k�5����N	�K󹩢X�s9/���I�G�&�&4����ܷG��ɼ߯��}�,MM����!҄��{lاT��+o���ۑ�9��}/�כ�<�"���d��I�6u_X�W���3�t�꺚L5�U:Mh�*{�L�Ug��� �T�-r �_k�y{��ah4��L/}|Vk�x����m�"��MTž^�^��8���x��Ӆ�&��.�}�_ ���}�bVҜ��3����P �
���psC�zn��	�����S�����nҚڂo�58|�~;�uB�8�3�����k��p��c�Z.x�:��E1�s�3!?�~����+JG��{��^h<1G�Y�6������;b� u�NՖ�UI!R�P��Y�B�dz.ڻ��XdZW�y�.�#9��&}h��S�$@��рub�_���Q���./�x��(�m��������	1�%*a+j����n#���I0�-$Jĺɳ�`a�&��n"H�L�����r�Yq�	\�=d�#!%�����t�j�oU���2��|�7�ꪎ�\,:����kI?n��nYx��з%o"��+�<Ҍ.�q��!	�[iѮ9 KN4�^�4з�}��a0�A ��zCHbj�{-k^3�������s|�8���R�yj!X����0X�;�����]��ؼM�	��hJ��	�k"�4n��~�$rV���eݡִ/���T��ID7��7�֨ݴ�ߘ��}(Q�R�����ٿ�\Wyƥa�ļΟK��nh6��v��3Z۹�
�Vh��R���T�u�o����$�񜏸f�!:G���E�:Eh�F��_�7�\!N������8���i��D��"�s9j�pdf�ק�Qǂ��l�VCρTl��Fȗ@��T��S6dPw ��^�6������3PmE�XY�)^Z��(����@oWѦ|��ɉ�O48�D���3���)q�C�;;%��̕��fk�ʤ�/���?�\M�5׸E��,�"�_8���{M�]
��(i��Q�n:�h\@�+�o8���.�&z0p´c�0�4��4�۾|n�Ԙ��p<ٓ����!}3E��(����OKP�O������K��b>ہ���RH/�t0��d
k�˭Ziҿ�D�Cٻb�&)���(s^�[�
���`��$=��+�7Pf�xb��k������l��J�T�I�h:��;�����l�|ٳ�t�P׀�p��c��Z)��|����j ȝE��yx� �����s�̓Q��ֱ��4�<
�^��~�E�{.�yz3/[�D��'fX��o	)#zF|�1����T�m��7 �U������vdfg<��x�#��%��j�Vߜ�=�[��[��q�+��`��}�e�a}���z���e�^�z���o?��n6�$�ȴ�����/������v�.�"�G ���X�be��|/z��͙"�?\�35`p# �F�4�!��Q��$>�Z+��';6cw�|��\�1�f�wR��Jc>Yt��N�����p�M��PQW�=��p:C_�L��wp?�\�Y�?#�*ؚV>�L�Qv"��ct{�S^҈E!q��ҩ���	,�
Vw���&3�cKEG�b���a6��H38{ߘ��f�#ͧ���ZjF�I��
�h�5��/D�' �GwQ��L�>^&>|`�H�]6�(�����d�n���f�����Ggڴ�w�Nۭ�jhO喬p+�K����o��l����/����+�=�@ ?*�坹�Ҟ�Q�I�:����8�Z�X��άH��{磬�IQ�� $���x:���G���n.%I�ɑ�B�.*zy�~=@\~��������Œ���{�����14������N< ��?��O�θ�Fh�(ڼk�o�C%����Aw}�?����^�M;t{}+�ǔn
Q�h{�[	�Gy[P��W�&����)�^QT!�w���ؙ�f^x�y�1��Vu��;L�˽[�l�"(�o���ʓ`�1�y ����;���h�Y�7̓�B��Ib��Ӓ9ǝF����Ǳ���]`A��iX��p�w�Q>�Iy/�	f�H�F�q�}oa�\@�f�r�J��RG-(�IJ�$c���/������6�@ؗY��8A��%:��M��g�;�:�,7o9i�"�;��^{�W[iIdǸ���;���jiH�{{���Xh�U��H�&�9!c@��࢓�E͏��tp�����Y���G'ۼ��Zi���؄JM��v��K��(���z���[9=g���̏����G1�*F^N�=}��yC[���J��
�
�>?�ws�\��)�|T��eWh��o��([4����ߔ���R��:��bZ�$�,7�X�
�7�E����V�_#�L\Y=��E�	��A��k�Q�}<J�4��½|@���A�}:<��3�:�n�)�Z Ctbn6L�m@ ��'}k�"+��4����S|\�l��>=ݤ���<i��cj�!9Sx�=l��W#sה��w��u�o'<�J!�,�_��I�$��o �X���q�G�L|a�4��֏��0ЅC��o-�aU�%��P�x��57���f�-K�s�Fsvv������AZX�(e�E��iĥ<Ҙ��T�*H������݅W��U�T`����Kg[�)[7G��>�P/9�I��K�6�*�?g�a����s*��7��!o��PxL�y��Yw�XI���^ݘ�� l%�Re��/{`�����]3�0݃.#�؅�q��_�x޺_��CH���)���F��~������i�C�Nfm@�Rj�PE�!��R��)��b]�lDoW�-;����q'ka������!}�������
�5�M�k�p�.�
1�c��3����c�x� ��C�z�`�_��7��²�u�gA1zTMZ��{@z��+�����1�d�OQ~�H��3�= a=sES[�R�{+���@
�90r�T1���o�;)�6�G'�ÖD�5�^���ۼ0�)Ӄ2��y���(_��1W�bƕ	S�(��6B���^�4i���ߐ��G�J�5[� �0����5[�$~�ڒ���������Xׂ�|'9(��)����&Г>�4�e_�Xvr̱��E�����>�r^�Y�3L*'j/R5��kJ�Dj����|K9B^���G�� �/��~����� iHb���WPy4��?~#V�o��'�shN��o5'��})��U��-W���������X�f��	Z��?�^H�)�}�����H�5Io��a�'��(����h��<��S�6:2[z�vc��Nt�)���O������o�X<�Ӹ�l�>�XWkEC!`�M!��щ�$Y,��4 ��+K&�#��[�R��s��(cm��?V%�L�&Cx�fzY�W*oeO��Tz^J �_��7]�*���ե��l1r�����Ȫ*v��8�D}�h챮u���L�����u�4F̔��EI�_집���K;[-[��h�X�vi������oD�0,$��|�f���B�d�����2�S[�h � G.#���Pf����!�h�ز_Q��"�|��]3��i�T D-~8&:Z	�����F�h5B�0�q_������eCB��>>=P�6y}O�zy�H0�W�)e���C��m��qɱb���o<���I6�;^�o#Y�ʝq��`��Il�=K"�r��@� ��R���$/tm�:��$�?��Ʃk���=�B3.����\�]A���#��⪲�ȮJz��V��!;�����'~o�^>n�����=Ar��U�-@a���>Bo���t�J��m��J"ݾ�I�Sg��f�;'�7�	K����R�(� �˦�q���.��*�U9?Ċ�S嗋��u`�}q/��x�n>�y�Q>�0�U�9�9�Wi3Ԧ;܃�F>
�v���Q[^v�A;ڃk��^�j��CН�=í�ꢈݥ��1�G���t��x���04&buJց	�}-��>��h�+?s�(�]Yݝ��=�S��j���w��tn�DR{�(C;D�$�1N{�L��Ђ�C�RL�<�m-�o%Q��[Y�?]1*��F�{�e��=HK��'�*��l9N�6�2�kidu�V&��ʙ�&/�^7�%�]��p����+�,����Q��|4(`�73��U�-�U�9VtI9kH6��衭�����,�a��R���G�v���^�*ne�U��	!x�<�����������_�hH�-�	�2�u��L:�V����<���k�|��xбk�D܎���h�?v�'X��󛏳�w��Ze}���S��� Sst yr��?{pB�˭��s��^�<K S��h�c�<nhS]�O�	��@��oc�<�"Ό@γ�硌Q"�2��o�����ϫ��8��6�.��*���� K3}�����U�8�7�ɓ�D4�A 	,���J��K��8�I���zp$�j�2�/�Bi�{�w�֑�N�&����PQ�unL��E��>�j2g�Fy�0y_S	�
��o܉�Y�2*��7�FLX ����;k2�N��w���y�05k�;	�XXC��}��`;>�v�m�i���ՏtJN����]8 ӝ���;i3s����C����ն�c�{(�u�#Z�9�Ҷ�쉶U��_�vU0��B�e����V����&r��G|�4�iY��[������J,���(���~h* ��@��޳�i:��?�ҒN�������B]x�w�3��x��j4*�Na�rV���pvگ7K|��:v���g��/��%=���Gޛ��y$T�n/������~���䵧��cɗ}=�t^��F�ɂ-XS�{��@�A�%�:��g��V�S舻T�5Lf�s���PJ�����&���^�>��-f��q vF j����oqX@��vk�%��Fn٤���L��_�;�Hc�啛&C5���!e8�J*�����McFAX���y�\P@�'������3"|f�J�0u�3ҀH��Q�A#�L���+->
�����@����\�a�����⤃�!��Wi��D�?�ýps�@���O	��sUV�%��X~1�8 ~��AFXgţb�q�/lq��w>��/��`��)075?���у�b~T��cS�~�5�箉�y��뀎7�"��]�=x�٥ܱd��Go���foP񆈰լbfgt��sc#g`��Kؕq�K�����p�}��y����j
p���Ч`*�]/��7�%��L��.R��N���3��C|y����I����g�~lC� 	nƧv��,|�ejް:by}���^�a����u�!�����U��Y@���a�#���C�.h'���&��:Æ�m�����.霳���2�c�/i+9���5�+�̳ 6�C`G��q	V�ꦊ�[�	}����ʛ<�}Y��3�F�X���=4&F�h_�`���E�v\('��zx�$"�qd�oR�FW�~6��S�Z���gxNJ�����y�d��k؍�T~�ċ/T�y�ɲ�T	�!Mu�.�3��ɰuY�/�L0Q��nK������,���4�UA�/g�eo�W�H�ߖ;C�Ǻ�\��S8��ԫp�Et�0�������u�7��Ln'jJXT�%����W7����f[nƓލYj����|}d"C��~1�ӛ�c�;q!�O�MЯ�7�1�J���ҭ�}-�r�v�Į�ܷ�!�J;�����iEU��z��Q��%<|66�}1�;�O8t�"��~c�/��
y�$�|%'���Л���)��!,?���ʋh�ģ�l�'k^#�Q�4�Sk�H�˳�׫�^.q'(�³/U!%>�=���_ 8W�x`4 ���o���)+�og���cu�M(��Gx�ʑ9'�������"{N���g�dr K�K�g����;W�� �t1P啚�&�fc�t�
\1�l�)�eScP��-'�f�(U%4��A�ad}�Tcf�}d�.9&̀, G�z9mǷ;ī�h'����4���C>�2�"�R��9l()�L.���5���vٝ�&'�!9�Y�AZS���]�s�^�	�;��u<���I�������e�j�y�!���m�!��`�6���G_h�ZZ޾��T��Q��x�
 V�ȯ%�J�ma.�@)��S?�r�Ȱ
!��u&�����,d�</1�m���G?%���%7n��k^"����������ˍݙ:��E��s��y]�A���9�]�r�AE5Իz���������A��)�9��qP�'~ 38עk�F$_��-mKH��M$�m,Y��IJ_�����D�Zw\>eFF?~YJ<o���S3Cw�a�� �WY6�4����[����˂p�5����*z�/D�!�B��K�
�rl0�)���-Ѥ�a{?�A������P6�V�@��6�ۭE�ң_Fz����6�� �5	4��4Gn j�j�ӊ���,"��;�f	..�Nӵ��2��%�\a�LJq��hʫ0���NK����H�RZI=F�GB�I	�����O5�%�g����3��+++�H��1Ju�9�3�D0�dZp�I��?�dՈ�g�����?������a�.�4^��W�R���ɱѽ����_�n�8h�C�Nɶ;��	I�X���I���-'�Q�� z]�E��]
{�Uɫĩ�B��½���w'��*+�\�9�ġg����,��k����׻��+��5�(~ �;��"ɬ�/{��󹜭�"�h�J��T`.���å5�	T�Ym�Ñ���Ⱥ�5鞞t
9fD�?�D�8�~e�1'0o����`�=������0[X'<%��?y%�F��L�-_���:|�*�{��#���R;{�f.n�EL�趽�"OE$s���'t�O��L��M,F���|�����O�|�6�^4vU���]oh�%����Sc��1�ߩ9��ok�<ש�H��e:T��}�O
��$eR�v?�lji� !n*H2s���eD�Z+d��QT����]=��O�j��_.�Ԏ�S���|΄�#�-��2�
�������	���>n�3��	����"�+'p�~S���)��(#x���l�.<��GI�2�5��.����IG�*������D$�K�Z�v��l�2�_|��K����$����m+Y%���UB�� wā;���$4�f����;&��L����y�Y]DmlFE7'9�+�Uy��Q5� ��z�T*7%1u�*P-���;W��-�4�~����nU%���Ǯ@�9��EV���$��U�[������
����c\�i3�ª�Ԫ�Bu1Go����ț�Ζ+G�G`^K���ς��*G̛�_���F�2��xw!���-d]�\��L��F����+�m�D"6S���N�rv3а�r.J�ڷ�Z$H$��L�礣2�)
FĶ�c��lv���K
1�d�N�؜R��e�j�7
Jf�W�G��`�s8��c°�T�N~��t��-/�i�����Z0ux1ӧI!��y<�
8�r酏>��H�R\�vвB���t�(�m��n�k�d����&�K�[�^����ȼ���K{�̇�tm�GPBg�~Cx�5���mWD*Gz:`���Ɛ��)n���IO��e�N-B̓�6�����h��Z��B䢫ϋ�Ng����KK?ڵ�	����QVjW%�~�	]>yCxL�'Ai�������$^���n!��a)ѫ-����5�+r��э�B�դD�^s���L=0�_�{}g�i&��s3S��Iq޷r��v���f����4(�0���1i�D��,��!b�b��n��},�V ��9K��v�|��e��'�����"c�
�x#���������8������H|�]q��Z���6��4����Dq���]N���g'��F�������\=��힡�c��Af���S��魴OZ5
������*ӥ�&*������������q�{�\mp/F5X��Ne�8�8F�]�^Op���0�'dX�M#fp�"�\5��~H��`�nt��U;Qi��'���g��@o��ש��˛�&ib��eմ��5V�c�I'Ȑ�u��X�Ux6�+��}xd�{�ï��{%ϕ$i{v�-d뚠��"�Y��ӣS,� 1�|��6ȸ�*�yõ���Td�Nw�Ls�
!�xX@��!����۩¬7�E�T���ٽ��i0�����pˆ!!z�	B�|��4ʘ~�J�������F�Y��ޤfGe!<���O{}y7�\1��e1r��:�P���F65�7��n$��ou����ҳ\�N��trjU�������6�bG��ȳu�����E����<����&��������R�ݛ{���?����������SA��d���
��CHD�[ ~v�=��>K��������ƪ�8o�4��c��eq���/�q��rj]��,�ъl!,�O�`E�Hp+^_��HM�G#(�[12���#���*�d���r�
J��	f	�"�x$�'�}�����y���N����hҘ˝�|Mq6���ײ�Ũ�獁q�*	[�7Ւ�FҮ��d�����*�|��@S�<�R��M��M���2>������G�E�u �o�]�������@
�Hi���s�#��v�{�T�T$��\]�I�祖'�m\�w�9�E^�K=_wa�ԕ�O�S~�(�Q�GB��+��V��ڏ"g��Y�cRX�Di�߻맰�P�uq�_�ݳ
&��/� -=�Y*=΁�)*N3~������3�%i��܅r5�8����%<������~���=����8A�u�w�w�Z�o�U�!g�|s���u���<d��p@n'�}F�*3��3|��R9z��4؎�X]ҩj�gF%���X'V��NR_��˕A��g5p���d�Qɞ�oJ��ݽ����h�ߡ��e�+�'��\=���z�Yr^�E/[��%�����N�|��W��-5�z��?�Ѯ%'lڐ��A븡׳��uq����&�˗c����@8i�a�{��!c���2j�K��)��4YH2�SL@�"��:@�&q;L��lTE�:e�6�/�X�dG8d�QV~�	�_�U=�]�~1�
2h@��'$�k��n3 �%#LK��=����\MX�v�T԰��F��RX���f�J�U�C��ӳ���[��[k,�V���F�Xtz���6��REe�{PcI��uX�2�BuQ��}u�'-��3��odS&lWS\��)_�f��Bl`.�}8;���Y �Cv@$��e��K��I�
�I� ᰹z��VƝH	8�bz �!p�G!"��g�(k��,8����4���>�V� �ݚyY=��^�=j��$2p��`<��]���X�*�V����$���#e�
�)]ף��W��v9x�C�w�k�f�@��C3��C�|�d��ZUǕ"�?^��D��?9[�:�8d��RD�}i�T�DR�OV�����ؖ�;B�j*
f2d�:�O����63�f��'E�����4��-����e�K��Ƅ�&�΍�����HžS'�O�z۲I}^ZO%��X6���tC�)`���A�1��P7����f���P���l�#���,f�Z������ ��u�TkGB��-�}�#�mE����1��Ï���°�fv�=Բ�^��Hh[�%^�[]�n��*�i�SDOP  &B{&�C*���x�p��{�k$:�d��3����X��&=�i_�('��k߭��PpԮ�ygiX�����Cn�j�"�"�[��
�� \�N��W�Q����H��*��I��u�;؄4��N@������9h��_J�j���|Q��X��N�K�!�[�J�Y�4ծ�,�%�o�-+��z��<��+=r[Ӄg=Ы�*7�'��SF�� �c؇��7d%I9��" ,��O''��c���@L�npI�fdV3�ݰR8&�� i�x��˭X%�,��'%�l6������zB^�|b}��n��c��0�G����{�
l�{�|6�<z�&ބr�=X��m�  �J�G��1X�#7��!�N�b\�eo���?�"(��������ok����r�=��ׁ�X� �����Uc�T/i:Lz����:ru���=��Z��HPBM|�U��~c����%P$���CT�n�Ф�l歠GS���d��@ұK▚�k��~L���-��D[O��6A��;�kr�t�d%3��d�����+�(yҷ���b��-�P+.�f
�8V�^z8��sp�X�T�A$��>��Ry�'3P��2��
Z�(�W?��Α4�eu:�%�=����27���ى�U�F����|L�J��5�
�@Vk�j�k��b$~޿�F�i��䯪䐮MJ��sB}�n ��w�Jf񱺓0_+��٣��B,�[n3r!vH��N��9n��I
^L�c�q
��h��?@R�z������E?�u�Y�;�t2)�RovO�>����E5�ΏT�
]PUf���0g������Ia>93�Ob<'����7z	��:0�M'"�� �<-��-Ւ����R���࠱8/"��۲� 64׻Y(�q�c9�Nڷ���虩�ј����E��'��q����� T�Z��[�d�(r�����hE8�L���K����p�N*6jZ�_���O^{���x	��gg'�^�JU[	��>���d@&�� �l*R�y=?zr�� ({o�tݍ��	l���V|�:7 �����
Оҥ�H��pƓ6�Q�dǛ�`�܂yPw�qf^fb��!��ckK��(�J���Y!LLx(;�~ݕ����b�23�/2���L���3�B���C~$4��1J��6ӤF�K���ΣZR�E���>�]r8熬%Uf2�g�˯��9��=	G����"�4���r~y�@�kl_�c$x�)s��{�@|��*�x�:��Z�Xq,.�CH�InW��_Ha���~����K3��uSP��/Ac�Y��9˅:coHh6�V"�d+/����p�[��"]�g?�)T����++k�o����8��Ly�,�t��)VEy_��ͯ��ڮP�v�j�,���W���5rg�ܙ��#��+Q����1{o�i^[�@WIa
@�ʕ��T�ζ%T��8� �񩺀���g��b�\N���Y;:J#\�
㯯���n=�D�����|�n��,g]����%�5�*�]��Y�R���)����G�\	k��܇�`��t��H�2�yه��E{�M������51���6*��_��E�z�	x��t�
���m�nښ�ِG�N�Zǜ�Q4�� `���Dm�O���QĜ?��a�o�`��b`���@7k�If����⨨[�ZVr�����܀˹�fD��=�֕_��E��.� ���H��2f)N{ߵSCD�q�`M�l�S��Ǯ���"dJ,J�,._(8�����P�V�:� �9��'X�{�.�TȐf�����J���%;���!�ĖF��)EvL{�����ַ�^��M��T�rk��E,N�VL�֫g���%� ���7&�ʂ�_�p]浑3�#o�2Odyn`E룮�[r�WT敨�#��O.Ex���|��6��6q&�u����雹�E���d(2��h�q,X��#tD�0�	�Fa����,�����Hw�s?���ec}��@��)��4��ߧߘ�y��}+�Ў&�+:@OY�wX3f��V�4X�����6�@�9j���;b`@� �m(3sZ��� �*�w��6��w-����z��U�����eZ�R��P����G{�����n�"�����}��'1�<Ɏ��J������^�yئMf���]�퐟3��	�:���|hՐMt��_ց�.�񊟐�>��"�@j�u+�K��}��$��P�DEYL��h;֢�N�w��X�ʭb��"�Q���`i\9���L�CA���E�O���d����ְ�T�[���Eg�Ҏ\�g'�[f���D��^�f0i\ �D,6g�'E�:ߛV2��Q��5�T�i[�S��+�x�
���-vZ����_��{{\1��$���xf���-�E[�H����Z����>���đm���I�p �~�LW{�w�}�+��-2�"ٌ�B�YW7C��Ҥ��0��\��dS�1g���c��lVE�nԗ�Q]�W�W���fe�8�� ��\ ����x1���}X<k�O�˒��m�����i]��G�3��66��&�]�H6�x0�Q��f	���P�p{-�-�&N�����?���D�d$$�0�o鳝�8�W�h����@=E�@�+M�����и|znx����K�+���C���;��|�sK[�[��e�/w���EDx�?��6�̦����!��Դ�]�`�x��(����pgAC�i��j��u�&�1S���vcx���}��_41CՀM�jk_D�B�՛��'("�bi���U_K��6���0^$��n4����EÈ��Q՗+й!�T�ՙ�gk!!�����;�c��6E49k��%p�Nߡ,����D �J�[���=�$��4�w����$ӷ	����� ���t�r��`,�Yw>�q֜���gqMV�x�A�-K��%k?�a����є�������ؽMI�b�_VY��. ��=!�0x��c:�@n�F+g��' 8���-q��J0]�ŐK+~��`[Zۅ3=�&8/�WE��&/	�9�O_n���!pc����m�G ;��3��,�՜7�U�,u�`�J#�1�������cC�yH����0�%ͫTKop�W��BX9�#+��zZ@��N�jNn��s�#PlT�*�Lqk2��|#j-�����s�X�R"4��B\ ��ya-羽nY�71�a�"]��������1= ~�+�Q�?�'x�2���I���/�i�V��f��SE�ވ���nCM)1�5%����3<�����Ag�j1�n�cb�*.ڗM��.�)���6˺Zd���[&�{+	���'��ݣD��8��/Z4e�Y��4���祐2��"������!�"�Q�l�C�!i�y�8��R��C�jD�x_y�O�'S��]�d�3����Wy�� g*v��=B1�^�ֳ��='2���7�f��"P�K��;0��U*g,��Ϡub�8t��2��Vh)իV�<X���6�es潴F���K�s�!��ɲ>�<�{n��7Gv�����9�F!��ȅIZ�I�P��*t�qȜ��G�g���h����[�\�1�Z��`u���/��h�Ӭ"����9.���l���Ǆ������h'�l�J�)���d��ݫ��=ś���U6��oP��m۞�������	_�dCl��;	Ε��|��p���s����Y8�Ȼ�Z�L���w�}m�I��9�BC�E�g7:��æ&����˖>w��˞���7�7��M?�J�х's�3���c��['rX))�y�R_8��T�MԉO04��fr/�O�/\����M?�}h��Qv���ŗ w/�x��&Z�y�(�6��?��o��H�"le!AGn���94�:~W�r���\#D:�Z�47}&7��خP��l4�S���)�T����c�䆕��a/�\u�jP�[�}[ ��S)K|�Lx�|�>o�^bL���P"#�W�ӗv)���� O5���ʉ�s��w�>?��HU}�T��^���U%�4���}s�t$V�?���L����,̈́ڕԪE)����{��n�b:�-��G�a�y�L ng0}O�\�v��Y����Yl��N&��x"3&��C�� /�%�HsC�*�E(!Ng��;�@�/ �am�����p�4k��n�^��#�p��W��<6	���$�|��T����Q�t�qr>푛�)m��}8I��}~�}� �V��: fauf�ͯ��S$j=M�cJ[���VW4�$?r{Ῑ�㦜=�T�`�����6�5}?/��!=�23v�%Ɓ�u�n
��,�� H�G�A�����а�d�/�K�5C�S��_��f���ܡŌ�ffb�B�d9�L(Z��'T�v~Ne��Tڦ��V�ƕ7�Ӝ��d�=����w��Knƞu�q�p��q#)��cQ���+���8	�}�@y�#��wY�2�����Ihղ���H�c�<l��Z���/հ!JD���Ynm1Jw��U�l
@�fɝ�jh`��!���yG������]����/̘��}c2$ӟ#��ɜa����Cj�
N��y�ҫ�a�j"|�ܰ�o�=�,��J���������o�*_po5��O�(�q�l޺v��"�WHP6 �)�����9���k��9���r�`���Y�c�T��&����wfC�^\ Z|%�O��Ѣ���&8����òNt}Xy�Fs�t���q��tKb$Z��q/쒀�m,��� z4�6a�p���E�C(.1���č��&�ީ��o0��X��8p�3v��2�a�J>)	��F��3�j�80e/}[x蟷E�>q'�\G�X�f����܈�4�|�s��!�c�@�&���2Qc���d!#�N�+�z��Q+e�_��u:�IZ��<�7O�ajҼe(��[  JK�����1~?=�j;�&<�'@Z���BI9��5�b�]$1�b{�b`<����O�R7�M����4�l�QЍ�(kry~B�����ƙ�=�E��"��|A�%,]Pè�5a��G�P����d>Ų>됀;��o1|�5D��T�"��B,�6ą�%l��w�Ǔ#�&�碫<ӽ����w:N��K�d:����ծ�\�����#�����*����d���~9��P(���D��	���͵��H����)B�v�
���K�H^,���\���~k0�93殷 �7�@�e���|��JI6`�����ٞ�9	@ωϫ��{8���+������������a+[�?=0K�Xf�>����y�?
ӆ�jbM�T^�B;��ʥ�*�Y�|�LԴM�*��P<�3-���n��Q6���'�b�kx{��'�[{�[�X�%�F���^�6OɅekN��l(���X��Y�8j'��&��#樂5U��P���즒3�1"^T�F�c�Y|G;��4����-�~R�0�~oG_��b��`2;&�MK("�a��
�0����a������c*�'څ�}���ا~(A.'P�eB���6?��4مO@��V�*H`���-q��q($�<��J��?��T:�޲�ͪVz������Q
o��0����,��}/��3���d�j.�} �<N�� �����Oso�`�)t�p���[Uj��Rdcp�ۡP��d��Њ:-��R�wad��ؕ������Z��V�$Mw���ʮ��+:���8�]��܂r o�箔6#�;����I�\�Mz�oB�_�:e0�~�����h�m�2�l,م���Ng
�)�?
+V�Q�r���1v<$A
�o�3&ȓ�52��Q`=�p�f�M� �2kk�󬨸�^�Y�����AâR�	����e�[-��G|��������ꐇKW~���� �/ѧ�!��
i��B��|�L-Rk)�|aߒ� �Va�0�R�"���[���������5��1�K�8�<��8��w�2���R�}�]pؤ�６c~����]M�81jr�w���
"WP��tH�;m���ovk �R`��ǿA~!su;��I�y��n5H����dU�T)��A���NA=��o����'b"Ǔ���D��:�zK��#�Hb�Oy�`��*���L�� R�6���q��{T�^�@x�W�XQ����K�ZrKl������ֺʶ�ī��s�ӟ���P�6,6 zb&>ӣ����/$���98o�r/���IC���M���6�2��~~y�C�eEd���ӝv�����7(�=��E�xA�D�Bgk��xαJ��w`��c��x��d�/�Tr���K5��`	/N4k�3N,���_�@�<�����Y�鮫���C���,�R�PӠw�ь��b�j-}"/G�;����I:�S�GR�Q������^�cz����\�2b�,ѫ�e3 פå�0,�Qrq�	&H�m'��l2Vz7m�-��J�ȑ�Ћ��[�Y��*I�Q���7�� ������|�|��"�M�Ѽ-� -8����E����S���G,W�,ģ�����ݔ0ә?˒�#�Ďh�ϕmVIA4�Ne�:˃�G1��_��=�Y�X��J��{�L�	E�Y�j��F'v�=��h ����w�-Ɖ0X�*�ӏ���m9�Ѡ=��Q\��N�Za�.H������m�*�5�]�W�\-��c��u����Yڃ�EV��7�x���e %�4K�/i����M0�ՆAό��V��ҳD�wsH�m/M2������A���	w�	�f�B�Zq�����rf,�ː�	Q�h ��4 �����fWtg�[��)�"?��=<�FU'�,z%�f^~k�@�K0����9A�C�i$�rV.K����z��{��K�	��� \i���Dg���!4����i�'�E�K�čխ��==�b8�|��1���^-m�[{�����h�
�̮��=�#���B ��:߽t<��`��D�iђ����1P��Dwh���\]�D�Y��X�{*��_@�k��5�\lqL�r���Rg�	�[�^TU��S�)(/�Qr�Z΍^2M�; �5lw����q�֜��އV�n�g����l���D�IV��Ԍ(�#���FN9�ő�>�m��nc�t��(ڰ@v<��K�	��/.�W�0��?�u�B(A�ŏ���h���q�­kNaؑ�W��)��2i�ݔjz`e'&���0ig/|Ƕr�5��ig��`�o�,>��j���J��[%z<(��)`J�\����-��X���<�+�ڛS0��6�E�㎿�ǫ���c�*�E�$�� >$Ѱ��������m���L���P����_Ԣ�d�f׮@�ͫnƼ�Ppӷ5��+o��hI�Q���s����.�m`�����8�@G�`�T$��'��JF�䡋`M���5�~B��d�p������Ĥ#Ƙ��0��z�j��6�?���=�k%ptf�ѥ�I�E�ufӑ�B-X���/?rcT �O�J2�xz=;�B%�u��!�G��k)*��0V������Zl��.�p�pv�{�'/g(ܛL\ž0�۸RҪ����R�{��3�`"�@�NN�Z����E�_M�[��$��Q�t���]���C	�� D�HT�Wi"�"�]«�j!�aǤ8i�n�X��Y<�΍L�F�5�1�7&+��=���ir0=�y�~����h}�Ի�,G�눃��l��*x�$�D�*V;K �إCs��f�3���$��9B���e��k�7~8zC[Y��(�i��2@+~��m(D*�"��r`o��Q�j��`
��c�A�EW->��%봷c�5��!9Y�7ѻ��Z��z�1nh�O���/#�ԕ��״GD��� �,�V֨�o��ۊ�c�ܞ6�8����}B鲇f���%�w�惁4>���F���`�d��0&��g*	�)��tC�S钬(	�=(~��Eo!p�\t <�*=�7� U�Ó�z#��9]k��3H4qmY7�G��琠_E�}8.>��SV>c�T�7<�-�䧎癓b���*�s��|폆��Cz���S;.���+��_C��gA�{�6�Y�Z1XN���g�/.O�:�dU��m�9��ϵoKnv{}��
N�r��e��{���M�jƧ���`r��/P�o;	@ׇR~{Y��[C��5�թ����z�f�F�\��	�rt
�� ��7��s�`�cG��Dz9��>��f�������,^u�E}`MJ��J��˚��5�! ^頴�u����w,f��KSGJc���� �NdW��\� J����ӷ��KPJ���v�%�����I��_g�1��g�r{H��0<��i�\N�,Zٿ�n#e #E2M��XC=|�Lċ�R9?nJ3�cp>��q����6��$"}����|d:^�
��r���A��*5�T"�I|��=�	e?A��Pw��Q��]	���g_d�Y��?ʛ�SgK��*8v���cc�NA�mM�����V�ǞC�1b��G|����գ���,�ȹ�5,ǰ�LrȽ�p���@��T���ugv�ݨ�l��In���=N�S��}[kVgydm`|��&}���rU{�Hլ�O��3��]%�rT�7@��u��3T��q���2n�քjx���l^0���=�	��3���qD��w/`E�{�6�<�4:�w��?+�j����P�sx&�R6p$���ܹ��
�W/#ą;�&�|�,��S�)����q���w���f=��$��,a ���xt&H���{*D�{{��ڦ�#�pa�R0<�4w����s�P�}xp��cw8;�]�4V���W�`阖?d��3F�YQ�j,��{��2�d��[9����K��`:�`F�%*IR�XD����+ՌS]�U���_�k32��s9-,��{��\wi/ߤ�%��b4��e��f�`���*o7�rA;�d4�.�Ge�(���K��^NF��!�^�I��P2̫}����7�D�w�P��q*���pf5#�5FQ�G��i�ꅼ5�zg#�z��xvQ��n�g$�`��E��z�v-<��Ǳ��FqEܨ#ksх����q���%���!
sD��obI/�Cԕ�S�� �w�t���y=G��
h��N��[V'��/
"�&?��Q�5�,��v�!Ta�o29��D��6I_��y�,~��=�+�Wj��N�D�橶M[�-O�f]"�������ݞ$�� N[�.}�!Y�uS��\��D5���1-۞uK��0\]��`����v�b ���a��ӹ�Y��!��?f7>a�F���y_�4`XZ)K�`3�=׋_#�̝3U
�iU��R �5�e���HX����is)<���o� ��y��fGЊ�w�3+���	i������������LxpXZ(���v����km��ŧ�,��f��q�����6UCK�8+g&��Q'�4uM�շe�}�F�4�P*�m g9�̨��6������Õq�C��3d[���'�f��]rFE{���O,���u��O��{��P%�e(=������3kg���c��?5p)�v�<D��$M,��n��V���ˋ@�E�\�S{�M�P@V�E40�đ[�����C5�f/�D�s��c�v�jT�4�j�u���'\#��"��x��)_�gk�L��2��N�������\.q�IL��NLz����6]����p�jّ&!\���ؽ���E����g�-�'V�S��f$��^������V�.v�'Z�@�i�%��P���L�T��rtw�nK�BP�KjT����Sԫ���Ņ=ߦ.�7Q'�^�;�(�hyF2m�i[�(:3/������S�z�'����FkX�Y��'�����d�X� �	2?O��yq�{����lkC �V�gg���ح*m|��nz[��_�%����&�4�p���])R�p	�E���"�� E6AD"k6��L��	ֱ�ú�n;�?���k���E��B#;⭖p�ބ*��[��e%�\����-u��x) A��߃E�.��*� V5��� ��D#��)9�IW���?��W���3��r���+��O[�w�_����\AE��8����d9�!�ywm8m�.��}R�7Պa)x;�����a�������I�"z�քV,�C;��B�lRjv�a����X�	��Bi?���y��L��j<���K�a8���al|jK14���x]B(����&v�^�ʯti��2����A�8� ���Nz�����ͬ���1�*�'h��j�4׌�����؋��pRǔ�8��<��Z�5x˴бDR�q��`�m߈t��n�p]w{x4Л@��P��-_e��esG�'�kp<؟6���7s?����vv�<���X
1���g�a����o�h�J���(��b4�J��o�k-uՃ��n��p@� ���/��,���a^�YuS�ܽ�G��>�#5d)��m�0��޳��8 �6��O�LRD�ڜ�m���bCƛn_���T=��E{GNUP����t#�t���ɳ��^+��DR�	�Ѩl9o)��Q�髜�%�F!,\��w��D�ï���Z{b]s]�ޝcA�0"���DU�����к�6�7��JƠԫ��ޡ�:�*u���-N!ۗ ᶬ�H �,zi����g�	�X�y�;�@f���uGSX�X��;]�~���3ft6�Z� �q-{T/NJ�3bq���CY�^�P."�:���=����I�����H�D��+=E>f@	����0�m:����k�Ö�`/.�������o"�YU���� �bx���-�,e>�Q�2��5��m���p��'jeQ=��?����8��v�\����|Sy(�
AG�00B�n�"ĝ?[�J ���$�lvVa_�xh�(^�{�\�$<�*���,�j��!�;�0)B�A�v��!m��8hZ�0B�������]�r�@(p�+Υ�q��V�EX:(�yw���nÏ�i�,���Q.!!@!ޭhlq퉗X�`�,�lE=�����/����褝��P3h�~��m�m��@$�-���_Z�u^������pM	] �92��Dβm	��`1{!V��z�|� ���Z#dF3�@g��!��# K��6�.��f�����ʔ�#��f�X�&�MНv��Rq�~���b��*��	���G
����vUJ}�L�L��4S�b<�����u�cx�������� �IV?z��=��Q����j[��*$(�q���F�ɡ��3��K�Z��+�e����W>3�Q�=����8�������P6�)p^\���m/�l���.����H�>_��"R��L��u��Q�Bs� �Ó뭫�~ Y�A8�P�
7�C��,u|h�� �(b+���B�����ɥ�����=���%*s��?i�]>��X�jAb_̞�`�>�mHEXE�h�9]�����2���C�D��S�L^"���L��w��c0HYFaq �\�ۧ2sB_S��Y��8RLM���K�'!��ғϳ�?���������Sz���*�"i��©�x�t�HvA
��$Ct�e�-�I�ͼ�yg5�ґ2	�x������F�0� g�Z8ϵ�i�e�>Q��#��-������(E;��;V��ه�<b=��ȩ#��_�}��d>y��㽉ƭ��w a,cmL���т���2�;���u�d�蟴�A;�E�����a/n%O/^v�[C�D-$D��o�9)�)�F+��
��|5�a�N�X;�ӯU5�I;�,�(�b��@2�nwS|�úz�>
��m`���L���W�"�Y�͠�z�Qs���N���{�yYmQ���₁ep�$�mV��YXʞ0!i}�������x!2N��~ �w`~E�w^��ш,�pW��՜��BF�E��<�]���6Qe�0oO.��Dn�4G�OGN��>AH�G���*V";��<�gb^8'����GЂ>�Mgs�ȓ3�:���g�/�>b����3�<�}�{q*֖ģ�U>z�>�jy��=Hg%�|�5&"e&@�wÐ�H�U' �܀������
Gxp�^�%�x��@m���Y���['�#�W#�#; s��F�y3�|�m|���Y�d�7�L�G�5��o}���@kB{��'g#���&;��nT@0�$&W��2�<.^���|�ze�v�5.�L@�<#p��3�=99�W�ȗu:��L�O/7q6K�\��p��ī��Q �N��f�HЦ����M��f@�ܝkʂ7���.��LBd�`����Հz�M�+ݳ��|U�	2��
JZ����H�6F2�j��|�����ƶP��$�]_t��m�qF����h�U���/�N������\!��"�=a����W�yX?�U�&���"ò7�b�7����[<��߯��(�����������Oh� ����D8d�!%�a�o[<�U��lh��R��(�I�ʵs��7�@~��`I�$;�Ocn�œ���H���C��]���1� �-Pl��I��I4�;�ڹ��]H�l�+��c�Z��NLDZ�灘���I��C�)_I�tR�YE�9C�)��w�A���9`=_n��g�<�%:%SdM�|���頔Ao�	����|��+��g�������N|�C�Gx�J�9�:���;�/ޕ�n��͗/f6 ~ӐȍjŅ�fI��� O�콽�δ+omV��T�8����;j8���3?�b���c�1.dߊ"��_]+��Y�V�Bm���ǌL����G]�q�_N�P==dX,����4m��*R|����N��(�L�\��Ӣ�OT.%u3��sl��9��-�?�N�����u��/!H-���3=i^H�%�X_�IP���1��q�7Y�`���{m8��mE��Iݿ�<1g��$ݫaO�.���ZUg9���c�Њ�-����È�͊2���C	�~�.�jȟ��j�����*����W!:��H���z�j>��!oM�bu��u_VZ���1I�3��F���R �9�n�:��v��c���tIODp��r�<k�������"4�� �vXQ�䠓_�����]��x��7��{���Jm�:mR�N��1ECk�����Us;mj��Vd�$�->)(�Շ�V7�>~����y��!Ք�����&�0�[Q�����5O��Y�p������PJP~톍�P�ν�^��ٕ�5}T�!:��ڵ�l���^mn�y�(2|���N���h	��Tfڑ��?8�D��}:��T��ӻN�JU�n:w�SW20���+3y��t$U(UAe��
i���B��r��{t�ݡ,_�� l*��[�d�0cxT$�]5��C��eÆ�1�����lQ_�sG�n�^�5�G�sF-�uE� (�N�g�,����{�ա���\�ƍDWܞdEt �K�ȍ�Ks�K�6�_
k�Ȗ[8��q�ƻ����@�Óo3�l�V��覗�N��G�+�Z�r��3��� ؠ�e��%����z	ќ{�*�U�7�7�Y�q�G�oPv�ɵO/�O���!�v������A�l�l]�уtw����锒?��������.G��d,hW�`�#Ccъ����^/����Rh��C�ܷ}�Z�׈	 ��(I�,�F����"l��ڌ����J��g ��3ƯVp�?x�M�~�����G �ο�^1��k9��^�p��oG�:H��d�@H���Jt��sS��~nM�<Bm�.B`|gb_7���e�Q���#�s��;z!���u��Y���;6�m���H�3pH�nGZ���3=��v&��u�w���?�C�D�B�T{�ާDJ~ܧ�t�����c��銱ҍz`;�� ���lgv�`��M���&�%/�W�q[�:��d���U�x�OV��;���/j�H�1%f'膄�)�3��z��1/4��1�M��R.�� r���|��� ����B�ڟ�-J��+�R7e�ᶬk|2_��R)gu����X�����	����(��y��X�h�;�v@>�J(�6�˜�J� ����y��V�yQ38n	��f���6oJ,.7<��xwn���&Ȅ`�q,��z:@����aW������{�,��|ڐZ��G��S~�l?~_�� ��A
=����Ռpxٌ�x��/�B��ݚ���S�����tT\��g&�)��)��t�@�vT���?����m͕w�A�̓���;�5�G,F������R�r!��n�i��Ŭ�t�	U]M
�<<�P�M����VD:�G�D�6�6AL.��������@�F�����������׿����5�5I����}Ռ��b	kD\����(V�e<U4�H�W�QH\�K+D��,�5����}!Q-��Ђ�G�*�Kѡf�ůt�ۮ�slTխ�,���m}5;+B��z��%Sۂ�,��y�RK���,G�!uߘ��^E�#/��!�=�:2�Xw9��<��Gˈ�]���i*\p.�vv�ٮ�7i�ҽ1t �����x<�[x<�R�J�{[rŮ�*�¯^:��s�R7^���61)PŉJ7%+�}�~R ⺐��TQ?_�}���Rſ�aM�y0��ʑ�K�מ�"���#4��n8�n�t{qy)�e��hĞ�A�B�Y(N+�\|3o�gtZP�s�L�>�Ę6�٤{B�d�sx+�� �}�̯�ս)����
�+�3\\l���3i�U>��&�ͩ��ЫQr�:�@؅BK��t��-�r���دG���ڌ�hN������ك�f f⣼R�ׂ�6÷�}��g���Ҽx�*a���g4ޅ��	�M�Yib6�r���v?�f�WH��p���Z�����w^��"��d��7��]Y��k��L�QH�?v/�X�1�^dF��4܌p0O�SM'�����:5�JFo<��9��ud��a���ܫ����sm����
�d�<�3��ې��g2���R4϶�lχFV�~�%%�|%��;�Y(�������=������Q7W�����'͓X�l*�b��#���ui�b�MDr��5q)w�E�H�R��C_
)E�S���|�����UL��?��;A{�$ҪK�#�RHoy"�v�0S�����(�{��\��ٯ$�����S��k�>�\�{}�?�`nbnHE���o٪��J��Yy�����j�;Ъ�)��A.ħ}��	��膔��l�^�֍c���ȫ�|���<A���ax�.οM�Ӄ}j�nzFŪ> �	U7T��Oif�@�@�'�	s�9��M���=����f�q!:��Z��/�d��>�a��#_��P�&�i(��Ia���2>S�@�v����q��]k�ׯ=Ϥu�!���,�9�Sެ��d<��^�<Ü,
���l���^cP}��}CY�v�H�ٿP)�J1#7V";����Rf�%3�#�9���b����tǫy�S���(�b��z<.��~��\d��u�7�������V�����Vt�m�32�f�W�"�f(�s�5�!��J�Ы��涃cmB��4�ـ���پt��W�3Ʌ3�=��~�8����~q�2�=X߁�%��9���͎�㡜���b�����p���b�&?��k�o��z-  �>lF��RV�n��4�PT�M1�S�a%k����W��� ZϜ��^|��I��J1P?��}+�nG��(���-��Z:_Ҿ=*�����&˰,�q����"Ogyf;,��Z�,�;|1�Ǯp�ζ��5�&k�G��2;�
4nF��B���:	Im�%5�npY ��Z4�sb�o\��NV�r�c2��6��S�s&RϻkT�;ח�VK�b���������[zGR_�L^L����_��'�T�ư�q��=����X�<*[Ȳ����TؐV
�M�L�1��  ��I�\����'��~�ڔ������?;���eF�˘���р�`�PDe4����%�)Z}jm�I�$8�!���l��$f��d~��L���l��z��i4iǈ�+�)Vؕ^uQKq
�vt8!�i�vU�_���WM�~�tv�P㽰�X(��共��5A�t��%[��^̫��"����B�)�p�*c�{�F��ULb',���8�6c�ӂk�ў#m������	�"0Q�D�X�7��}-��=������~���q辬�U	w��ϩ� �6��[�;X���Vcm�5f�ٮS�M/gf�*��H��\�ʴ+��D��ҮH�:sݚ̗|�o19�p��b[Lb�$�`�I�d����>L<�ߺ:�fT��#��lD!3y�9��bf3br\!Ӽ�L��Oh��[�N�T/��
@� D���J�ZӝvNf���8�u	sP�LI'a�SW�_#F}�H���ѝ%�+��'x��in�6�6���6
=+�&ݘe��[����2s�:�']�&�8g����©�T���ϥ�����c-��$[�B����P���QK=��>�9���*h�Ҭ�,�?������9ACt� x�}�<c7��*��tOp*�[����%i>e�KZb�?��g�B֝�"��`� X��R1���>%Cgy	��\��_h� �sD�<�,	|��>:��Eױ�G�t֮�(ޟI,�v��B����xS?�<����uT%	{��4n��B)�v3�hR^)���ݧp��`�e���<�$���]�*b��(խ$c4��׫�u���Wǎ��55<���T��"�Z�@h|�h ,�-��R�l�
�ADw_��P�$�SJ`��#����Y�a,p_��u�E�@0����1�����F�;�A�2/�/(���H�6��3�kꭅ�f�!
���p�p�fgOW�.��7	��p��g�3�Y�g�fZ��Q�b{V.��J:&�0�Ug�֍�g68�Y����+D�h����Xb�n���{��є��H櫏���N3��g5�r�lL��k�ƍ~�F߀NRΛ2������z�:����cب �=�$p}�����	嵄�����C�:��敟�,_���7�5��ˀ�D��÷Y��<5�����y\�����#�N���<����d��:�G�.Y�=���Z1�{u�.��-�2FY������W�D6=�fY��|�  h�	Q��B�q�C�0۵]�?��lR(;������mw��q���_)��a��R����Ve��h鍲f�v]`0��'��W�6pn�\А�3%ӆl�R9~g�>�S��^�|�Pn�\��n?ZBl~V!�6>=��(.�͟�-:��I�BR�/�8y�"��uQ
��)�n	2�i��4��#f�\?�XuB|�@D�#�+/_
+e�U%��M�3��$b�>a�e��4j���n&�{��L���(/��~
��Bև=a-��Zo����mp䀍���i{t%��g��	��?��e4���^B9��D����(�5��o����}��y���&�{��F��Nr���嗰�'��!�	#+�j�E�̞�����Ke|�P�X��Q^�a�ϱ��(�Ze_�x��X&�&��8$�e��z��C;��D�qrzO� Wb�Ӱut��l�]��	�n�}���ai�m�/��8:�<eu�9��l�E¥A���@zf�����6K��	�ʄi�d=�s|b��Q�Gb�5Ǐ�?D�"ik٭�d5�L D7Ŭ)[�9!=@"�u��$������,�yKux2��jG�M�ARw틼v�Y�ؚ��Bi��M�]N�;�Q�6�R��J�s]Z�U��B�lq����	��b��&��P�Fggi��L]D�f��2��R�W���a�&�݅"Qux#�q�׳%�f�Ua�K���,t1!���)�T�PĮ��zVš��KiJ�p3�.��t�r��H�%A	?�ix�̋8Ѐc�ECS�7M�094��g�\[vd��eX涨U�jG:y*��GP�nS���)�%ޟ&3�Vy��JFn�;E\��y����@AU$⨄��P�!m5Q�~fĕY.�<*��uui�?6��v�Q�W=2���M;#�Y�&P[Smw�<:;\���y|<�L	#�	��$(e�NR���"�ZM)� �N/,��h;�#Y[��&Q9>��j��5�ق��IV2�=C$����x�,���q[�>�����kܭ0s,'�C	q�kNu�OL)��K��&�����y�S�����aX�M�q��j�!MN�is�ۍO�\/\D2�&kj���#�O=�L맶�IU�� ��[�U̖z�1/fKW��}����.5;�D/_:C�(}kh��RӣS��`��7���y��N5��m������2/>�ߔ�2y�#���M�����E�Ej����BO_�D�ty@��/�s���~��:\�ɗA� \7|�A��e8�/�Y�^������5B�M.��Omn>��©��Y����01����f��q��b���S+J��tI����v%wo��A��L�"�?��'���H=�*���4jj�`����D�7�{,"��֜<k�c�I�J�����ڥ�6��G,�T�H$��"`���B �C�敬���`�؀�NmO�2�j�ǔG�dB�M��3s��Ux?�8Ѝ�5+V������P�̬�k�:����A��S�l0)�,�ly!��`�@���f�GL�Ⓙ��j.n��?���>F�������^RkZ��˘�9�)����o�n̿b��[X��m��)c����N���H��2[�P6�G�o@Jnd�-����[Ɇ��n�_�j���x1S�7��j~�(A	��O2��J�'�G�c��j*g�:��_/>��a�$/Z�L^\OY�iR��+��:}��b��5*$������^�t�?���1��&6�3�B��`�3���u�6d�H*��̎���4s��L���N�� Z���f ��rS!>B\�=%I�\�U=���Aw�l���sM�+vd::fKw�s=��˖�P�Hi}QS�F�ӛS)���աَ]�s<X�g��~��	d���i��$�J�]���1�J�`�^>����|z��Y{�F�R����g$��9mI!�,�D����S"g!tq΀�ߤ�Ay�W�H}Δ���h?�����
0*i��Ҫ�1\�@��kΡm�m4�܀��L|�Ng�a�B��m꿂t�o�R�ߚ�40r�2Zĕ�h(�%LB��PK���"IGxH�v��ݎ�Xhw�7���*#��&����c����O� �l�z��͒T����H�V_I�f�7�`'�O���w5d����#M؎m=}"W����@�xm$b�#���f������;o����olf�$�-�v��׫��X��^�|4�q�k����GAkI?Ëu��N�p��X�!V��-�W��gd���d�63(�Rґ�:��A,��kb��v�}������r$�,���OuD����"4�N8�wu]���$M�)��������-�[�����Y���s���^�AX��kK�,q5|��a|]MDd��m��Z��%�ӊ�K�y<']d�.
�[�&��y�E �N���Z�����[Ӛ��{���h��k�V�e��`v�͑<:���)1�_x�U�g�_ul��ۨ�E뀬߇�H{�����΀�8g�";1!�b�,*�� �
ȭa1k$�o��"���|��9�p,�
?���_��@���e�����J :&u��a���R�񒾣���S��[5'�|;�)�)k���|��
��+{�� �d����l��P���;�S�8��#�
ǧeeZ���Sz��4L��75���u�>,�.-�t���;��S�7�x
��?}���=s���2�{s���p"RX)  ��s�����tg��(	b����.���
t��G�D���������(Od��ؠ�I
����z��W��g� D�,�6W��h��N�{ Z5.f�b=��g3�yhZX������G\ͼW��	O�^���Ѷ�gM�8�/�w�\��������c@OɮV*�>�4��V?i��P��`�odmP�#��?^zVD���t�*������z��B��T5/�ʻ��b#.��fs����F�`�{Q��V���"Y�<���ARDC������\�}.��4�Ƈ��d�>�m�,�������[�H�!�p��?���'ؖ��*B��:/gO�a��ل�0�(�:7�Zfb�.�/�����)������֔��ɸ{sr�L�b	|sc�R�Jg�h@V��n����OofA[��o�sə�.�F5�G�G��i�bXye��/�H<��D���1U,���жE�{�����.U�=�2�T���IR�HW9�y��HG�T3�)����`�8�L�ѯY�ld�H|���ۿG�#X�3�(r����`M������j��a� 1�P%�z�ؑ��+��/�Rk5���nc�t�6�^Y���$���G?ʽS!24z<Os���i~S]2|0���y��N��ڬ�K���%��A���X
Ѿ��`����@��r*߳~j;ȗ{w	#?=�-'���[�6��E��pΪC��>�Ms�V�Q�i��� [���K%��R�dy�m�F5HH�~��F^"�/§�U��Ӵ�����(&fެ.7lYE�cҦ���X���J�> C����\҅b9Re�2��-k|�_ ���//�K)? ԯ7�������Y߮��ȍ�I�2���1vP�Y��9����?4e!D�=V�3#M�	~�6_�"��3�����全)6�V���l��m��v���p����8����փwW�3�5_M��;-}f��7Ԟ�h�'�ר�����`J��]ȧV�����r��m��R		k��Q�:��3��I��@z5��k�Y�u��Ø�D���=*Gű̇N�p^�d�W���#�.n�)Sa��D��]
��"'�*9��'��J�M��&�M`:��5 �)Q�i6[XKx}�2����1�bmX̼����DP�56��wސ��|q֒ꅻ@�VQ���ڴ֞�$�i�a*��5�f+뙊=H^''l��. ��7w`$ϑ-���>�]5�&"�ND!��i�Y��jk'7mU��Ļ�Sy?J�X�+9e5i�P�X3�b���Q�M��܌~Ń�exFt�aU{�D��>�e/��o�x׷�jyu�z���������m��L!L@��?RBd��p�.g��p2=�hc���HH��oIs/����Y���fͩ��'��������ʁv}L��N!��e�x�� �C��-<�4��|�V�5���xAx(@3�8Ƀ�ًdy�}�R�fNZ����z[0s���p{�u.I`���O��hFi��
��^��	#��.�d!��
 ��1\�����`+~�; F�0	�AhT�F�1G�U�B��`)���Mqf�O��q=��.w�S���JU׺z'N�/�<��W�&Y�-�!������\�=w,T�&՛��jp�G�
�ڂ/���D�\�v�*��Q4�H�o��u�姱A({�Z<+�WVDxh2`���$[N���pfSVA���������2�ԅ���;�����(��A���B����1_v�O鮥��zM�5/E��V]̆'-��^W�����"�+�������Q�qz��B'��BK��|]T,'�t_yFq��ji½���$��f��X��g��Q%=q����Qe��1�6�UR��qXA�fTB�0`�>�}�x~�-ka�T�M��5�ڎ2�W�m���0�W�9yQK�v+h�	�����S��	��!�h�[1W��#w�j��j鉮h��*x��cDd��������������ʢ�k���'��u��3�Z��_Жm��9���U��"
�mj���6i�2\���NcE��>���U�9�F���N
%�/�Le(�sb-�H�_���H�鑡ϑ��W�P�]��%�����a�W��%�0��'#�m��G&7w�G��x�e��\�!�]ɖt]�G�*B�:��(�F�`�Tn��#̭��.�}�A�Vvk�0өgD*���5��ጊ�f�?�^��kOxtO�<N�&m�*��@!�{�T�7�z�=��̹�&J
'Кn�V�Ľ�{כ9u!�VS��a	�ac�5�+uX��ݖ��'�oD`�������)�t=�a<<JP������~#���c����O��$P�;��D��!N�l����H���g"����v�t�
[��D�3V�A���jWێ�DC�9������>T܅��ZP��'1�%�s�oB��Q%��Q���D\u]H��n������A�٢y������\���U�����u�EW6�,NE����G�ZI��Wq=��r^����_s娨̇�vW�}:����2�Y��R﷪���4+s�����]89�-�H�j�uT'�fm�q��nq�҄���О�r��.��(F�����&����8������t>Н��u�>|����t+*bt��0���vA������`"�7��>FR�Ye^3V7([�'B5�m�>P�;��u��Ct��������$m3O}�U�L���>%�nr,�~�4>Fm��WU���Ţ�Ko���%B���6��,�k�~�a��)�5=�·<~����3xc��'�I@rG#�F����о]6����V�z��1W�G�չz�v�I�_8�i�� �P�C>���eG/~�Μ�t�]$7n<S����<3hP&�[�cAtD㟷�.r��F���}zҘ�|��U��d�U;��=@Q,~��U���A����d�V���ɄJ���&�H�B`WfF͎m�Z[�ZQ���헄K�'�
��@G�l;9Z��@?�ք���-��(��vZ|G��N�0SvzO�H���D1cM�g��ꙮ.��K���t�2U֑��@�Xj�&��i���l��c��l��\�5B=��W3>(����[I���a��)��>U��T$������*��.8 S��QֵIkv����:.�P��@e����Fӯle�l��͝k��0����ݶž:�P]L���!��і\�J�s"����'�P)2�%��\��[��0��ZL�gv�:�V��{�	a	S��<�_���e�ZR޺,cwf�8��;M���y���s��;����C�h�ͧ�w�G[�`^p~30E���&���z�W��B�]%}ȿc+�?v�7a���[a0H���ſe�{��jŵV�L6��ٗ���ɾU��ſ,qຩ���,���3
u����M�~��;�k�����a9�Hi�5���#�4;��}��b��~���c����d�MAC�s�9h�Awprc��|�cop���C�xUd�����Zl���mçfs�qޮI*<ł�o	�z
�n:ꤞ�U�{�:	��T+P��G���Fo��ʌ���>����=��8T�w���V���)�XR7�9U��X���ߵ��d~�t�.��(-�AH�,"1�a��Ѯ}y�k�b?�,�����e�z��˕������6�Y���������ġ�m�t4M��5��5G�WD[���M�l��;}��� )�-�4�4��.����\ؠ���]�����C�?]%�d�l${}g�ݴC�H�ʑ�rm8�L�w��%�_��쌮�o�.�����v�ԛ�i�}����O�b����\͂����'�ս�<_V N�����_�c��琞�#��>�����'�#�JU+�����sP�o2pw���޻��"%�A?��x�}�{LV�Hh5��-�d���:Y*�	c�U+%�[��Հ?1WX�V/D}���o��N������!�u�E���{niT����E����|#��ꀘ��%�r�Y���7�Y���W�3#Ф���V��J�����i$��5�~���
 `R�ߊ����d�}'���¯S��п� ��*�k�I�%� ]������LÎ��7��ߓ葻�b54����$`� ;�u��,%X��~K�E�mG�u8���#t�5!U����F��bez�Y�c ͏Ɇ��N͵*͟�'A�Ñ�T|�h�y��2B02Io�-z��LiX�� ��vV�._"�ק�*nD�5�B��j�h�/�/{7���؜f�鱢Q.n�ziv�	�6�z�s"e���բ�j�!������=.6�E���R�׭魑����y=¨#d��>|s�cA3��.���^�;�x�kAǃ�'_ٽos��~�?�4+�V		(� �v��G�~�S��iy���ÆJ�Q5����3R��؅ݑ�CT�/ƓM����3|�"1��� Q���g��"����wGьH��~�Z? ;3����J+���ǶX�f0��oӥ���Ğ,���/u��Q��u~�n�%xe�Y�b���,����7��Ĉc(8��ƒ��]�c�NP���&��P��|OS������?(�x_�,L�k�tw鮜͋�6s�l���\��&�����g�z�%�U�Y����Ս�|�uDbE5H`�ME�GX:�р�:N�̦��,�K�
qز-;�W��>�[��?�e� ��	כ��wT�|���a�~@'���#��	��F��T'\5�Ep_�æ�@q6E)�N	Ig�b��	�t�\�������uV9ަ�~l[\�w�wd4ϖwb�ϑ��Y���Sm�׵���b��U8&ħ[ �Ϯ�z<���G81��+�1Rvvh��oX<`$��*���-��Z,Ҋ�����S�]���V�|'?�!fm��y��Y�C��o��o��S��B>�W&���ݶ�+pN�6 0��w��n�����������&��~~*�dn�"�mU��S�2 �Q�����5�9wU�,�lS�϶%�H�OG��zR��ۚ��i��-J���I��IC��1¢�	����ė��AF�p����s54v#�C]Q��@��j�y['���*S��*�����*t�FQ����;Eײ8>�7x���6��Dͪ)b���e�r��HԬ�D�����g��,֠�"���Qw���`*�[�d���t� �x8$=a��Bkl����)�����X��PW�؄B�d� �~K=��m{M�U)��r&p���k�n�-f^$LW������J��/�5G��>WtЁ��ey���}!�L���0�P��Ҙ�:�l��0C1zeh�%�Nʞ9dj	J����W���u&i��oޞ1�FR��;χ���[���Ol+be05�@��`G;>w���!�Oa���,!e����*n׶��R&��I���Pb�E�IȱUl�A�@��UeC�~h���;���Մ�͊7��	��Û�~D%������	����yߦ�	�Ϙ�)�#�,j�i~q8���Nޫ��<x�������_Y�J�=2w�j&���Y%��3FH���<���}�3	a_�wO��l�W�pj�1���Ӿ������(w��A�����q)��@���B(�K{���S)�˧Y��S�%WtדƼ�rƝ�P_���&9��9�R
�Ԡ�P�17���M�K�&G}�d%�iF
UT�X�lN̩.-D�N�#��I �'L4�U*Mș��`	�[?E�>�cD��F��ьA�@��ģ�ta=��ժ�{[���z�H9f��IX�U�8m3h|N����?kC���R��M 'Y�v��~�_�:��{@uB�`'� ���_W��|Ib#�f3y2�����P=T5��6^����Ƿ��˾�t\�r��i�`P��!,.���ft�d��(>���j}'}���I��?o�|���k!_ �:.�v�Ը5�2y�(�-x6TL/�&�:��v�y�v��Ne)���-a��Ϋ0��-s����J.W�e�v 6�i�����q@�7L4�D�gE�iȲ$�(@q����͌�mW��C��VYV���aҋ�g�SKPb�O4�<�ݠ�T9�z�pW秨��=����.�؂u��d'\ĵ��Z�<��M��v#�W#����V�W!A�/�x�D?W�T��=����`#�3��KT�Hk����q��k����D�vˋ��a�2�o�����J����LL�^
�j��&��M���s5u9c�!��L2���_�8�(��6i��8;{�l�%�փ+s�n�|T�`�c���O1%D�b��ùJD�pٕϞ�#���j���ֺ�\1�����JP�hi+�5sݎQ��Ev��+�<ݚ�"��_��r��'OC)dmz�8*�f0�r�l~��Ԟ�\:b��1�@%�;��ɟ1����G�=rX��q��tN��#��͚^Ͷ�H�:�O�	�D�c@�U+Kr�]\z �[0��6�\����_����F$����Σ4.����1Q|a��q:Z��OԪ?`�[�g�{���q� /��6�Ө�Ԑ��3��Υ�Z�(� �ַ���L4=���o���������r�3An�Ml���vo��HA�{����'7���K���S"]=�G:-Ȣ55�/%��՗"?�8�G�`��'����z�p�KDh����� Ool<���tMw49b��k�r�Q7IӀ���ܾ��y�YϠ]���;ʐ�@T�:k|j�O�Sک�ZdTn�ݖ�6�,��Զ��U]7`Ga�l��J���e=���0�ݹ�[W'~e�̓x碢A�Ւ�ﹾ�7��f�Cqho�R�����d<��5h���sqw��K�Am�­�z���31�Ȋq�-GG��d'V�El�`wF]� ;1�S��K-f�wox��VYM+�ȸ��RE�	��6�yJsF�s�O>P/�����A�˧����/��@mO3� ��u��B1F%n�6/�
���*s:��q��h��c�J�`�4�"Ȓ4.��/C�[���������k�AJ;�^�:��9�Se�pf��9�;Y�S��='/���7���'X����s�H��Q߮������:��탮���R��6�
o��%�qU��Jjb�-/�r��|�����uE�#��7�7M���\��m��oC4���QJu�*��FG"C~PzwV��k��]��;0��Ie�B�Fx6
I����I ��b��C�)c���n`e(��U�o�ҟ���k��2I�jI��7���@$�[|o�=5i�f`�m�97�
	��Ž�M�+���s�wj��רu+�4s5���T���J��MDC="��x-R�����d�gnx�:�X(���#ԃݥ�^ET ��j\R+��9�D�W�E�3.@s8g� �4�Ҽ�����q��3�ooY�DƩH����3x@��r�����/O���R�$=lٺT4�˳��)9���tK������{�O[�������:���+=����F8�}��*��<0�҃�S��m{3]��C[Us�ڇ.^/jRM���d�=���z{�l�n��}zK������thwOD0(��\���� zyx�7���!n,i��I,8?��'�䃕5�����p��%`m�?>q*�q8͐��_�^����B�i% �l?xY��)���� �ܣM-c���f�� �a�~�\M,0r�E*F�X� Ss��ٝx2�g�c+���E9��A�Ak��ֲjR��ӥ����7����؞���Ǟ�FH�ga�G��1��>.9nu�z� uP@��m���H��at�X�,�t�lMC��d����6��| �OB����� ��f2�H5�X�TK��{�Jx�R�X@��i��s,8X<ꌸ� �գ�U��V���o�69V:`��Jq��x^@l��2�n��V�Za��m���� {���$�Le��W:��1�n�'�e�`�{� p�,�B���F��o�ռ)�/zC���=g�~���Ӌ��s�5�72�ܲ�oʆP*��q��4:�V���7�JrTH��6l�g���0g�� 46���C�gjq���;�{uk��{!�ʅ��,�i�����AW�,��T�W]�@q=��G:� �#*@f+�H�Q��_�3�L�z�}�@�?�qP��������W�
�:#-'*gGb&6ң!U�l�Gr�x�w�nhV~7h��}K�p8��a�Xw�ߴ6ȑ�ַ���R�.���g=�h����"}���K�X�G8*+�d�F(2��O�OU���E�	�寗��˾:�4�A�5��L9?$��	t���o=���V�S���73�]��{��^�
�$Je��l��f:�J�1i4��=;�7�����o�V��`�R:o�"ɲ��H?�lp0VdH4�r23gV�~3���J �ڑ�d&e�B�9O5�+��I�\U�s~�Z "v�A�Ax��=.iuIA�8k)'�w�&b)zhGǻ1��[��EO;�-$A���BGf���
]�!��߈�ϵ1`c��x'��m(�����e���r&���;�� N�C'=�Z���k,��UU}����U����u����"����0Z�3�����ܤP�L�q S��N�K�ҟ����K;;YOMF��Ŋ4IͬV��>�̿_h�;����w,�&w8��H��+B|�,�)ka���"�>8w� �c<	w� Bz	�Ή3�%��y��r`@}����K{-$%�g��*�5n����fL^ky9r!�ܼ8Cަ�,$x��<�����a�пz�i>W���7Wւ�%���#$�n8�A�[t�mĕځ�|yf�Y��_����E��6�c��"��И���P&����9^=$blf��ǟ*P��x���I�
��Q!b�*��F��Xl�Ҙ�+��u����8�
����}@k��M:�_��mz�<C��d�^�Zj�^5v� ���'�����r�r��.:W��	�4�I����Dd�m
ԏ��į�&���������s��9�!{��k�~ww���a�G�{���ϟ�cH+�(��и�� �@������T�\�R���M��Ϙ��z��&H6����1K����:)S|�p�N뀷�����Q�)�0���ȟ�Xjl��e���z����31&�P������i�gI�Bȳ��~E�93���-땘�u�H�i�Xí�vy5��8�<��i���K��[��a�f ��(�z��ѯ5��:
���|�8a�';{�֥�������A.k����v�z�J�p��',!�̫)b#֤,��ɺRŢ|;�c���9I	�+��Rg�v��e�007:@���14��i�k�lm�cxsÜj��d:c��:U�z���ӷ�0���?E��B��"�Z횕�IGe3!߅��۳�@�Q/~��i)P��Rf4 ;�PFޕ�1b����l���ă���3:�T"N�)�$n�����]S\s�{xq�Ba������w�e��b���\�mkb�[B��PB��T�&��f���Oh�P�=�?�e�e��)��ICCx�`}kg�����K3�g���ߟ�k)�+eĘ�yH���g�+��s~����bM��8?�w��j��*��-LLBe��ͨ�ZP��M�.]}p�
Ք5�i;�?"���:�ܗ�:�/(���/�<S������l��L�<kkZ�m�m������M�2ڃ�q��-M'����d
z;k��1��u�%K=
�3��<�ބ�$rH�"h�w�i@�'~��w�6
�A�A|�-���&~�p��|S�i�Q��~�hF��Wa�d���W�Lh� "���[��~#f��">�����H��g�꒺q���n%��f��ۑZ��jhǣ(�$/�Tmd�����$y��'�@�����
	�O�\Ruu�
�P���f���x8>�Ͻ��F$z�zLhH[_����� �6QH�ͼ�D#�h~e8�-!�'���SV���"p�^1���Ft-+��q�h_7.��{�"'���N�Ҋ�8��t�vѭӰ��T���6b�,����BP�����q�*�Fx�����yT�A�e���r�|؞�+$P��Y�BM��PF��d}NQ�b��W#�ˇ�"P,Ź��>!x��%�p����N9c�L��^�|���z�㛫��x!�^;��KFj�6��U~O�����.�#Ө��u�*��堈�׬���;��3��w�17V~^VTKJ�_q���x8*�|���Oq����ĝ���WT�����o�_64�J}q�	�A;t#b�C�#�%dBd48YH^Q���F7�NYLE�yx�VB�GU����P�V�����v1�9o��m����.1�,��߆fZ^�;�H펻X��8Ԋ$A�!�E}g2z���������-xRH�F����m_�߭�C�)�p^V4�p^�/�`�,���b�UyN�p�ј?�[x#����Va6
lZ1UI�w5�W��[�W3���O	_���!�8^}�H�s��	���.�}'�uq�KF��^W;��0z��R��S̤e68p,p�<�&k~�Ȱ�4}�u-����3c�� ��s�xont��0w	�8��{V�֝�?].5��lK�k�z��G�'a�r�����nc'��UF�+Y1�c��nT�����}����m�����-��(c)6-mnd�	U��9Z�V�H�~����Q��S{�>�R�':ԫ@=�[X�y�Tq��4CN>ˌ��K�v�. ���C�yΤ~�)jt0�W8u����E��[���l�L���Ɏ-VW�Aē�]Ȃ��7�'�F�d�/��>7�3 ������Me7���zOrl���f��1��(A���>�=e}5	�֡�L��%����N�J��__��K�ߵ�vn"����j�AJΣ��bZ�����S�=�����藳rT)(�����\oH��8���\����DK��R�B��na�"�@���Hp'�R6B#�����0�8�]�${f�s���>Vn�PDu&�y�R>�:��	�{z''�
�}U�Lf�BK�d�2M�эS����?�o�\�LN�/?�����:f�pp5��v�Ǖ\e���Z��HӜ�D�L�p���̨PV"h���ᝣ�b�z��X�v�˵��b�B�z�}p��Ds"����m�#誈����9��$R �
���6a�`޼��6�l�r�t����%�,���\�iBAF�m��$&4'�6V�P�J4M�*�(����H%2Vd��x8��ѽ�f�&�c��r�ch0���E��J�@�	�tw���'��A��&Q�hX��;9��,vn� {�[���U*�@��)�%�0��
*`�X�bG ��f7kFd�Vzc�'N�e��.�P�%s��ַsT�? .*u��z��Ϳө/�>��ӥ}��
ɮ"X����=ڒ*��b%����n�Mg@����?"�t�zyq! {f�#TK� c���Ȧ��*x$�G�/֦�`a/qk# ^਑8�
�6"/�b���$��8���Y�U�RοQ�93W1KJ���	|��
E�k�_�by��%,�B�t�7�v��\sRG_&w|��B&Y_&���9�-%7�\L/8_j��Y����5{o�����#��T���m�Ish0�}3�E�kyJ����%��g���Ǧš������K��Y݆]G*h�i2^�bXM�}�o��Α_����a�?w�$jӿN��f�)6��.�����sI��d��L��� 06v���^�#�]U0|�W Ei�}Q|e���G�W��%��A��a� Be�۠�u��`R���$�L�Q?���u���E��2��(����v�S��Ωj
u�&��ǪAʈ̭��4��nfK�ܞ���2�r����׎}��ƺ͇�4��Cf��q-_8_~U�����%�7��{w8����� �uP�٫t/ش�t���m����rx*
��RTb�v���\>����J��v���u�{nR����4��	��7��.zxz��XI����D�J�[d;�-�$P��h����%'�͸R`��=7��R����bO<��S�?X�%w�V[n�j�6;�aJ��`��n��r�\2�=T�D��E��8 �S���y�: �xp��ؼ���^�px�g,�j[�P���1d@����)	h.ꁾU�k�-����� �|p>myrl�~��أ�ԋ~aJ��.۔$q?���jCp��`���OZ-�VӒ׷`_v�7K��E$&������a�}_�!�Ϛ9���I,���^�c�խ��C�\��Z��5��q0�������>1Sl]&��UV����`k��&%�߃y�)��j�۹J�>�̻G�3#W*yh\	�w�_Q鄪s&�.�g�@.m �O��Tc��R�9���Ԧ�;��5H1!
N��4fWB�v��,5��޷�c|�?F�(�CUb�b���Z�2�E�%Wsr%oU��i�A)��E����j��}s-Ej��,�ߕ8�{1�*Ҋ�\	��b0�>��Ԑ
jr���V�ڽ�]�Sj�
gUQ|;�4�*�D�ƹ."��g�a��z� ��E'N$SA�����Cy�=@���(�ƈ�2����Yp�Z1�ۈ��"��g��3��N��ITJM�-��;�	�������-?�$clPa�XӾ*s�|��Q���8֌���30a�iVk���X���������DPǳ3y�b���������ݟ`U���i�c��R��'��� �������-��*SR�vy�J��� ����lI��r�����g���pdb�TG�W!�ۑ��!�ݻx�%<m)�  d�:ހ�o��ǒ*It1k�/��,�C��z.�;	�#��i[p4Ҿ[��?�0�vj��x)(�.	r�7�1�BU#Z>`K	����=��/��b���Ȁ���?ӈ���A���+��%A.:L�?�)P���?��[��!T���\�/�������"�� ���6�r����A���"~�sj���.d,�7y,}^I�� �����7nx�ެ��y���F�u�Zx�����l#9����P�n���\}�QX���M[�sw���ܻ`T�Mzv>��*nO��K�����*��B���p2-]��ӅKTH�>�/ xv-�t)����?,|Q׶0w:�[�S��ţ��è�Z\9U|zj�(&��/9d詁B�M%لxfvk�=��ޤy��`9�o	}��MP�_��pS�(`]���n�M^e��n�O�q�� ���>�d�A*�/E3;Ń��0�z��dd�<�=���o�8~���59pȕr]ĸu�ƽ�$UNQۧr�%�,QD��p������^��Vp~�)zmnEY�$_�v���ȡBtV��`����"��:!�4�Za}�i�̬ G��<p�&����5P�	RS����&��;���ی�� h_ֹ}Q���b�y���vP�U�oᛙFu$� �)s�oa�������F>bp9���z� ���,�%꿝��mpϯ�t��7�di��yM|%��?�l�H� ����X~��&
�~�_,:��x�J����8bNs��y`6D�6��m�p@j,s١�w�亰�ֿ��s��	%��ŭ��::4��� D^#	���an����<	�P��-?�6:���bhs��5�t@�6������y�b��X�uMfnU�u���:�a/=g�~2R~��3��#�3�_Co� ��i#���a���ٍK����Z��<���b�u��XI�a���@����ɇ�\�do$��G�����|�;1䄢L��:��[}�<xS��ұ��%�!"湎� ^2 �SC��Ld������}�l����s��yί?N��av-��� ���LV���)�k"Ͻ���O�e8�+J^I��f�'��d�d�l=J��6�|^~��Ѓ��x�6��C���X����~S'��MEۤ~h�!��y>����g�.(��0)����Q�`��:���a�F�]�8k�%k4���B����y{��?�e]+x�?��w�=� �@M�	Рz0��W�t�&�����~����/��B"�w�����B̬:/u^���_�zhȌ{(Vإ��z|!N�I��3����nk#��R$�*�Pf����~�}�9x�)MO�	>���O]�d���h���(%���U��7�O�k$i�#}���Z�.�^��D"��̪��;�5�)a�CIs��4<fGpc���)}�S	Y>���꾖mM��t_ZK]��U���\@�"e�����ܝ��mQȥS����� ���]��7E!P�|���U�>���qõ S���\����2�"�!X�I)K���>:�y�]h&��q�=80(�p�*����F�T����n�n���z��ǰ�e�A��Va�B�ܜ����qӧA��������i^���C���pBQ/�墳-!�j��п��)���e�c���XH�\*�uE��Gh�>�d�լ�a�!��2K�58�|csY�).<*���;f'��(��n4)}w׿Q�w����̱9A�-�������؜X��W�>bG^��c�]6��J[v�ӌéACqG����b�n+g�T�5f��3*�,����uA��)���6M���.z����XEn݇���]K���բRsҳ���ZU���֍�:���nU�`����|�K��yb81vy���d�s����Wq�!-~��R�L@ŕ�� �Y��_�Yc{��Cd�`�^׋2��Ӏx�nG��^J�SS2���-�E��r$�$(r�RjL��t7`��b'��݀�U�4/� �n��;���܊�S�+u\V��g��BD�*��O'�*b�Ԇ��h��X�N�CH���<:WI��f������9��n�f3�M������Վ�)�Z_�.�t�  �ɳ|Զ��ڦ -W"��tp�l����X:���8��&��������d5!G!�0O�J��Z�%-V��|��o|x�-��@oI����6�dR�!��L�}�5�� �!܇�Α�
q	�L���>���k^X.;u���N%z�'�����e�mtI�W�n��}d��g�d�|�6y.VG��G�8ܹlb[�VK���h���{�K���@������B�f������� �V�\�2u���;K����gh�������4QJWpg�Ȏ_��=�=e.0�;L���}��V��ka���0��M��@�HQ���D���N�fж�9��*�ۇ�� ������:QL�|>Jk��B�\X��S$A˜��}:�'.<&�
�HG������8V(����1��"|HH;�ɣLQ�Ұ�M�n0QB�&݁�-3�J��E���視|���W�"CA��ذ���9J�/M��F��X��̐
�'1��9�*������X��{|�p�y����,2��k�'J�Fi�n����Q J#�9iSrܔ��Cv�K�3�� �la�w��\�B�y��?����)���	.�TkM�N��Jh�N"cc�D˷��S��Z7�|�����~���F�S���Z��g��_jb��e�����=�bV�fs����އ?S_������1�U�
x�I�U'b�)<'6��#�J����m,��W���`��`������̢j/��vT���6-E���ܡ����i�D_��k\���x0�Ę#�\3�I����޼
���+��nz����F��H���7�� �l+
�u�m�ҶN������L�[���X8F �ɓ��/R��Y�(�k�W_��*��v���d�,3�t�%�˄�D �pD�5�k�fO����Y��*D��Eٞ_��ˤ����DwpC����p�sd8�X}l,�6ń����|���>�6���ρf83H�FF(׸:d�0:�\�g�-L�9�����wl���K���_P�I��ϔ�G�S:Ü� ��7��9����M�� ��u���m��:bq��G��e[TD�mV�7?N��"�b�6r0s�J���`|�%��L���[T3BV�3j��1�:���HMr"�	#Q��������մ�	��;F �6D$@���y=� J����M'���������@`�^�%�{��t�T��{6&m�2�d�+U~�-v����D#�j�mw�v-�E�w���G�-8:QnV���d锽�r��K.�m��%�����a<Ȥ�pd�V9}��n���v�K�D�aæ����K���~�iӺm������ حJؔ��W��Z��\�3T!��p�������=Z�G�r
�����=��y5�xa-Z�#��ڧ����ԦVe��.���̾Z���urU�,G�����V�z�ՠ��K'���._aZ;�1��#<�WN`>�:�u�1M�UpX48Ʉ�1=VR���l&��Y��E0@��r��*�o{q�+躺�u�3��"퇫�D��Y�� �ǁ=�e~
|�>?B��6ݙ�%lg�~��O/ A�qU@� 7�7��mCҠt�����L����ΪT�yY� vo�b�/��	[��q|N>3�$7|�2��o�qg�4ֲQf>&Ǜ�ZJ��O�L�U(R���h�O��SXk��*�u��K��?5�7&N�D�S+����$/RL��Z�(�@F?��:��:��nj �`b ͌0�̹Z��̥���1�}�� �l�e��#���j��t���68�d@�����p��R]wIW{�bj�-���o�k��z]����O
���C��f��:���[��dZowI�|�iQø���x��v��� �Qi4'�&��'�hWz&�P�";��Oj�cN����
����v~�X<,���^�P)v�;-�L7vu���Hd�F�i�l �:f��ԤD/iF���VżPX�ᚵH'�Q,���{�yd����>����I�#(|H��Ub���8�s�In��})WC1��;��MȤ/R���:8{̺�j
����R���m�]��~�9��"��3�55��3hk���#k�&Z���*���׺��Ar���X`B"�I;����!+�8K�0�H�!��"n��O�od]��@/9j�
��tؚK7�2�vY�',�&�4j��Z��4�/J��p�{�U���ڮTK�O��sǫr�O��"��Q(B���IV����t�r$�%�t޿�,10u�5�������j]	=[��B�X�<��Xyҥpm-�Q���NU�Byl����?{Q2�|�=@P����慇X2�պ�D$���(���w�(B��`�ra��Y�s��1A����>*��
�o�0gwd��b2.�l9��_���٩�_�G��(��v{�Ԡ���/�Ax�PL�$�D��~�i��L��D���9��<�pb�*��3#1������f��i mwz'�h�>� Il��X��b&wҏU���No�6L�E�\k��PY!�n�s-�0<����/�+X��\|hH(�eqF�w`78 ݲz����X��8K��Bɰ�|/w
)���a���X7�6`ko:xSfh x�4��o���bA-�y�W����rة)�^�2b����Ѳh��LϹ���V�Be_4�|_9���}X�4W^:�l��H��.�$�I�QR�~8R��<XZ����5�4so8W�8�[IP8��2d��Sl�EA��g�����Э������U7Ptz�Z5"Lĺ&�������`����B�B2�yl���ll���I����s�.I<�q -�K�������(��A�IgC���ެ��T�A�s<���s�NT�����\^�UV_�(��E��]�⮎?7^,��1��lP�R{�Pz����ݖ�F�����X|�bBo�������5�]�؃ՄkOC�qI7�D���x�<] ��dx%�{G2MT�L�E��AAY��AzK\���$�몿zka'!2,颛�&�$|C�ᅙ��6�&�p�|r�ʑg�|�ؒo򢇅j]��H�D�����zt��CR��Ge��]:�3ɳm	�;5�ċ�s&%�0D����gq�,�G�\����qytߣ�<^��CP�0���p�?6go�Q�Y����W4�أ!����dgL,�u���c���]$�|���3�𝰇Ūl}�������tt86H�=}�
�N(y>���i�8��*N����^�@	�D7�Eo2n���S}��k+��ߧv��V�f���m�s�O����VYV*����Q�O)~�oh�ƻ.T4��gG�A,�H鬥�)f��2�'9�j��r��|j�ؑ��a.B?�qvQ�v$��6�L�� ����5_S�[O�)�Y�4`���n��j��ked���n��ӣ�yDպ�%ѠH�l���8�6�Y_�;>^"!N��b.~xA/�!h&�u^Jd�Z��D�h��TϦn���j@w�uqN�	�\L�8<�������dʠ\>ĒO��4Y�-�ΨYM��d���Ng�d�L픳}�%m��g'����X*o�V؀1y�6%lWQd�#�e#`��)���/9Ԕ�F�+�b�g��<A��W���L(wQ��1�Y�\Ї�gfFT�
�����4�V��p��#�?�P� ,�a�P�_�����8��1�S'wK:�� np�b�Jg�����Ec�.�#�%4%�]tz`ܙcS-��XpX�p kV�� -��Z�b�H�jnˀ�_�`��VT&7dz	�c�~a�3>��	�I������lj"Csj��)"F�[�]rr�ʩ��~��qs�pQx.Brg��^�G��G���cXM7ǖ�T�,�)�tPd�YkA!�Ɲeفr��*x<��!���B�y7#A��O�Rɕ�N�P�J �[#�d�4"c�W#�9'�Pɱ��Q椎����K_��D~�Dϑ��i7ѻ��}�Q��#J�M1�V��Ǩ��a�7!q������̓�!������@��09�rz�b�p��&:e��ϕ�P�Z��0��H����a�\o"k��c|��Y����z9*���(�5ܬ�I%�e�Ur��, ]��v���:Ͱ����"�2�e�j!c�]�cE�T^�+n��A�b@r�3әp+�@4�@檺sh�s���<�U�l���3 b��3A�N�,���2�1� r�'�xh��а��޲q���|U�N:,HXYY��W�<��M2B��G�Jߊ�1v��.=�u9�t��7D�~�'fslX��`kb�t�k3q�Cņ�n%ٛ��ʗ��r���c��?�o���~�$�}��w᝭���tS��yx"��jH[��j*��s,љG'��o����xsqӺ$�^5|Z��n;{*�8��2���J0�*=0"�엳 Z��ccqT��`�~���s<�~�])�2Il9�$��Q��{����zQŒT]A��jL�m�z>�������B#R�@u,�:��W�߷[��12I* C},ў����r���,���;a,�*}$���;��)�J�-㾨��}�f�0�Œ�s'�:�93w��4>!�3�ʅ��u}�OgsLMZ��-�t'��dyr�����
×�P�r�G��od�U����B-J'2�h��g�����;%dL,	����w)S�t�U3
^⸳�D�2���|>��w�Q6�	&�FR�O+�̱J堧Pa����L����A楥�S+G�Q�n�|2��$�j����Sr�J�&o�7o8;16��x���e�Tܞ
��M9n����0=/IH&�`��"�1i{mJ4qϢʆ��u�V'K�;�j](� ��rg�et9^%�J�g�Cp��տ��BӚ�6wC��gЭ�z�W�+�M�S7i���D���f���1�CE͓'����0�-�D���F��P�̋!�hR�!u����� �(T�V6��r5i�T�J��=�@�β!h2U@?�7�x��E{�1��)���^�5$� �����8�A��cԔ���<2��s�a�i�Ttn��fN�=�3����K���H/�=�ոޓ�#&q^+H�,M&�&<��+��V`�o���\���P9����f�%����-	��PE���+�m����k��O����g�χQ=�)?�ȑv�%�b{m�����3'|�ˏ_R���֭�;<��IH�E]��Ks�� 8D�7����+�{(�HB�u˕��9@�v��Yl,�nw;݋6��;��]5kƀ0m���S��G��u"�
�$pb��f�	�Y5��~Y��+ݵv�$��u
bZ�X@������c���ɹ
 )�=pjO�� ��|�������F�hD��3O��U��LCy�!��%�K�j� 4�gӾ��X����*�~�$��=Ć%��^u���u ;;�Q/��;�l*)#��<ęj݂x���Z��>��	�YQ�3z�����S̶���{lV=`��O~q9�'�zk���`� 6)��cv�6d��󡛾�x��#1���&�������=�:C�$�K �`H�>c2H[hz��X1D���h����§Ɋ4;�A�\V��e(�q���KQ&h��Z�U3���sٙ&��R&��$��ȗ��_0Lur��'�4DR����mC&S�p�l�3��?!_�nA�)u��O��oe�^<^Z���b���T^$�D�����!�����i�)h[��e�?d�m����N�B{Z�D(���%��k�����A�p=�f��hX�t�[�\������X	����ɐ<�j���T�����:���e��T����}UA���X@9F�W��!�,���ĸ���yE���e�J�![�H�i�{o��Jo����1Ej�˔�fr�0 ��=��	b5��^8�*Y��N�[����T�oF,Jt���� ,Q���(-�c�Sv�]���� 5P-Cb1P�ь�/Z�&��|	m �� e���Ron�q�949ȩԮ���Aq�� ?��r �,��g�;�,�qy9��*Ѭ����}��5��+��� O�R�s0�>A�X�}�Yk�3k&��5Fk�ߎ޲k�
[� �e�i����s(j�C�}V�����}U�Xg.�������bvb�w}wO)o�"�k� �F7e��YWnu,PY��R܉v�w��U�,M[dm������N� ����nUZ�@^~�/A��U��E7�qO��{�#��_r�#�$ԕ��Y�U�xRh�s�a�6u'4ZD�Q%:E�)��F��ZZɌ�x�k�r]2�?�!l]�KV�	��l=e�AMC���CA��<�
���%��g�d��"��Pli?�<AVx�KW4��u�zb!3���6j�X���>��7%�7��zJ��c[�FG�ؘ�cI��{�a�|�V����x����	�(�9ɡt�����-�d���?��a	����W!�15�]�މ���J6x��{�L��co�O��1C��'(�v��8���B����I�	������P���E�U7�{,���j��Z||YJڈC���8>�s������!s�ڑ�Yy�;�	��; `�^��k*j��߾���)̤��@�L��ē{ -+E��.��TJ��m;̟̈��:P<Y�?�J���3f,b�p�8u�T�g�d0퍂~d���-�Y���L^���%��J$]�I+��溍�j���
�UtT��W^����VD1�yqo��i�?���7÷U�{"��3�r��Z>����0{/ŭ�s;>��
�L�X����|�1,�����������\���2�%g<.������rT��?�S�o{5��]�oMH2�	���ilm�!��\�Iw2��~4��5OO]�n��z$�d�+��b(�#�Y�<�i�%���-���s��Ϸ�����,(�=o����fFR^��\��g
OH�2��pN�i��H���������m�7�nR��~A6�g�<��z�t'�&�>K�lG�0(�f:bf��e4���<h���߿csG.g�]�j��GSd�_����H�_vև�-��զD�3���%�	+W��W��?��b�!_:>�9����v��f�n5,	(t�X3G�G0��M��ԽkO�OhH4ȕ�7A�֢-�XL�תYeř�Z.�����xӱzT䨚�!�]�V6���y���C��I�*��Z��j����9���R�A_�R�3�,���p��?�jo^��+W�K,:�O�5�w�?c�[�L�sp�k�e�����_�~�O~�V5v�Ɣ����/�:9
|�c�M�h#V?�Ύ6_��-@��q�E(��B�~��Զ��8����|bl����g�m�.wJ3�����!���a�)
T��|U+;j�\}е���L�e�O_a87�i��b�Sj�NHr����i�#PeXM�T0� �Q21T�B^�q���Ѓ� ��Rzg���G��h�!s��Ϩa�]��̱��ja��xj"�~�Ĭ��*�@����S��9����1V����ac��U\�A!��#�Z�Hw�ˌ�#�,��o|��۶�\{YZ��ls�ps{��J��4�4���7H�h����	��랼��qz;,�\C{��1ĥ��}錪��ހ�՘�ߜPݸ�:ꅼز�;�xO��.3
V*�$�b��P'�1�H&��B��7�hK�A_T�Fi�1��~.�#��2����Ҟ`zYs(mQ�j�V�+5l'��^C �����+2�����Z-$˻�k����K�4_e����y|%h�s���o�W��q<TP���[%sB��Mϟ$0�T�����#�����K�������t����y2RYh����^��m3v��@����svGy��J55��Ci&R�����Q�b��l��o�996�2���78B�� ����uo=���G��V���D$*�F�a��#r��V6Ќs/��Hp���?D�Z\>�3S+��`�����d��֬�Lk`�7?�������`1��MiO=Ql`����9�V����k>_��èU"G.	�n�ݷ'ȅ^C�[�fN��d�_C���̚�Eh-��y��<����Y�ʄ(��F������mK4]=��}+���I��(r c�
�W��u�^nr��2w V�&�"5���Yh6ʥԘa��6;̻���K�G{�7�s�3�}q)�b�-�<�>��z{�*���������"��Z}>xs��"��8��*Z }U�����G��F���M����u��@i�%��-F�0�_ڞd��?������^ט��$;Go?]��ҳ�������^z󂷽nj#�[kP���^��B��J��Uk�N���<������X�;��5{�5�z>���>��_j�Zmb_S",ӌ�1m��8��#D*�ZߚX��FQ���<x�R���_�z����ڒCY����~>������m�]�n���3��6�5���~�q��+$��A��2?�G��h��B2I��g˒����v�C�'���	��ދjo��>af�X�f�cXD�:t����D��P|�&N��^���^��B.V7�K��$������ȀBB����
e2*�.Dk�H0z�>+lBx����"�GP����@�D��<K̛�+��	��AD̫���34{e��z�t��Y�o��TS�D�DX��� ���sU��^�A�1P>�1S�D�ЪP���&O�o�Q�}nM0_�q<wy�n�(�r_��HXt����;-F��$����lg��� �`�@Iu�SV9A�<����՘Z9/�0��B�i���F���|�]�v�LOfuv|d���#Yf����֐#9v��p]7vi�����D��泈�S��ǔcޖ��E2#XS�XV�[�5�o��d�e;9��Bأ���M�)j�Mf׿r�����K@��4T8b�4jp�@���ơ����d�v�	�w���w�?����(EO�$s9���0�	�B-��jt�*F
��:��l7~Hz�/Q�{!�kx�\<7�(�{ �R� I���K%��$�b��,E��$�|B~�U�([�kg�����]��j���c>��fEƵ��'%����ʈOV��;n�:+X��^MR�����ډ �TX���b1Cg�������걬:2?��2���3@�G�`�&�@������ �틵+^�w=s����DL>��2�~����ٯw�����`&;���!�Rݰ��f���nn���H�I�,M	LW�8 োQ�fO�����S������*��z��P5��/�ҽ�K78��f ��2''�#�ުx���yD7�.�͐�+��� q�-������>���&��*J��5,�SV���~K"zZ0�{z9Uܿ����mM��$�0*&Z=F�$g�����"�����Ұ,����]'�>=����1�ǧ]:���	����
��̣�К������-���|s�Tp�'O�1�	�\�ԫ�~����)�Q�Lg��Z��z秊;����"�>�k��n/Ko
f~]�Oz�����ρ�ݣn�WY�>�UB�LPi�*~��g'��������_�0�L��i���Po�y�D)l@�Fؙ#�-����qGY�ޚ�}$O��1^�|Oz�.�;��Nڶ��Jjb�m�vzSW�ou���O��02o&x�љ^GW�^f�f���.�������,SɩHnT�D�Q#�Bk�
�O�4<�r���7h�����AЈgt����H�2��#��V%��t��(T�t�C����
��'�{c�	��u��T���	҂�N)u�zW>M�aoF�6�v,��^�f�a� O��Y�2�ӌ6T��_��IS_�LI�L8������T�^��O9��v�*�}6��ן}&Y��0��:x��N�W�G�ԭ�jyM��k U�	|P������o�7"�r�!��N$�`ޮ�!�����,X�{ڙ��}F�s9,�~ ���I��`����"�+�)������$��wCT��\�j��kU.�E\�=|2�He�ZjZ���v���٦T&�d��/��?M0o��O�I�k�� 
��d�ң��զwǒ�z~�W�s�o�6O����R�nDЧ�%l��.�x��x��l)V9�+�y��T�㰃�C������٩c�w�_\�U}��#�_:�GI���uc�*�g�%%�uW��$8�ct��Nϙq�I�T�K�J��x�%h�<Ԫ�|k��h�Ji��ry����i��k �1�I� 0�F�� ��������PW�s��Ŏr�/+/�W51U�Ȱ�_�ޔ(�]�N�x�N��|��a�]R)��;�胡��;��ȋ�ª��B�x��i�/���#�cʦ`�p-�8��c��x�^X��uʧ8�^���P�&��:�b)��Hu?)�;q�&�^@�zY�����`��kӎ�(�gJmsN�����=�~4��M
��@;LVc)�:+O��ׇ]�l�Z$���G`����"� ��ƴ���\��P�e�c��ios���WPo"yL4���X���zұ��.�M���ᛞv�t�y���/g�M�eo	���M+^c�$m�b䧚�c�#:�\$e���t6`��=�5�����޾�*�6A8	��^�:;�1��$��q3��1��=��z˴D��n Yw��Ľ��1q�ءV�%�������wȸ��\�y�>���P_�./%���G�4Zm�)! ��#R����\�,�Ǹ�ZsnH��{ph���V��Ǥ��\jP�g���ͼ�T���x���b�/�D���0��Ўag��86�ϑq�Z�~:L�H��l�Ŀ��Oø�I�]j��6�k)��X5��*��"H�X`B4,y�t�Ӑ��f��r��)���� L�D(=�B�g�A�����W*���Xx���i�O���i��Z��43�Û���) �j���wK����u_�U�=7���C��Z���\i@��͞y���Q�UD�؟< @hC��GrS�m�DҘ|@��  3�n����W���=^aPhk )Due���,���=u�����]J���I�|`�jo���[u��Ϣ�7�0���x�������D��&`>4�Ë(�4T��.QNH�i$��ّp��G��d<*����7ŷx��� ��2���B�y�w�j�IQHԲ����~��5��}S-�8p�2�1?,j�+�ٌNk�)�Ѥ6[)��N
�5,�3q}�5���(�)�h���T��<+�4��y�C�������k���UE�v��0B��X����-k�Yrۊp{9�0(m����s뀸r��W��/;��#�����Uh-�_g�,a��tu�{�:.^��r,��X-�:!�2����%w:��k��&!�`m'T8 c��0�ԙ����ѭm��d}��Q'�x����# A5/����6_�)Q��vw��gAg�g�T������o�f\Z� ���6'���$o���{;]���	/'��?QN����<3ȶ�MF��|qi���[�ȡ��"��Z������PJ	�Z㋰��ĺ���]��Ic�S�?ʺ���+e�9�bA(-���t.�28�{�%nk�p?l�R=�n-d��z=;G�#��c{�BK�����L���M�6'lɠ�B48������>��:X�4��FK|�B�X�)s��%��}/X'=Ý��K���R��	tN8I��ӝR�\�
=ө���w�Ϲ�qd&�,�TN�bC쯦�������hW��Zip\Jt�w����o]����ЭIZ��mډ�iB*��\XÚ���Oac���.�T�MjZ⬢ywf�\T
��I����yq��G�����$w�B�!��~j���B�dQ������Pn]ю��U&�XS�|Y<�^�tw^��v��IЩ��2@4E�����>8Zل����PYKWIX"z�lP� Q?�2W���\�!��|��I���BG'̇�"O{&7ȝy��b�h���*��w�UBp7�8��-k%��m9пw�p����z��qi����C$�8��֏�ʈ��ħ�Y�w�f����(�2�|q�!�ae�h�����[e|��H#�������
,�X>,� �N����-2�Bᒚ�=���>����L�����f>�%~ݾ��$���1��N�L�Y0Eac��y}��C�����X����A�2���9�I�	U�8�Yg�!���c�&��J��d{T�ݱ��t�B%TB����Jg������5E;GUWR�d.��4i�La®2����s�9�_�}	��7�:.�?�aE�(�Z���} =���?���a��P����5��n��3�|�������r.�	�]�w���~M.�W8s'�6�<��0���AF}��k+�8��&�ǩW�f!����P�c2�&�ϼ���H�v5x^� c�>��58�g1�$9�59�U��y ��wҨ��>�>��ӈ�x{�g.�F��W`A�Ej
�Q��JH��r�(�Z�@�OQ�����@~<���Y�RblNZ,D�*��v��/N��b3n�D�1+�?�\-͸�ǝ�NSX��
xYD���v�y\w��$`F�l�V�Q��Y�h҇8+���������:P  `��*J���VtԦ�*�L�������A�9�L�����D�F�F`�T8�ޗhe�-�ʿ��Oo�_O^��J\_��q*�991��$�.NGb�X��ʊ�3�#�\fU?6l��0��!��1���3��~xr?6ʪ#<!����|��[�^���̷|TCHĉ����LВh�S��Z����m�M,�S{3`ώ���@f�#QH%�*T#( ���J��QB`4=���z�Wy@���K��Ǭ�}��s�������KCH`�T��S�z��d@~�f���(�󼑡�������H��GM��ކz���I��z3Y��+k�MI&+3Sv�K�^�&��}/��	E��D�D&X�qAQRM��}�5�вEt�Jt,�*��娣"'Tʱ&��`P�p��l;I�=8-���:\uc��i��KĚrX��WX<=��Heq8du��&�d����R��+�QCSĈ'��}��VY���p��8���12\�A|�����P���'�����d+a�zh �������qXBͳy�6�_ٶ~��=(���%�5V�m�������u6`b��F����Oƌ�G�"H����4Lm��x�U?,��57����s3l:@�O��r�Mx��'���b��c��<Z�����5r�T׃Ed!����A*q�X0��{�y�m?PAY+)�`�\�����ߗ�<m�v�g�[�~���M���j�؈ŗ"4��=�qq���4p��@�ʱl7M�k_��!�"�͈�cb�u��5;Ov�蟂�5=� 6��Ckf�3�r9.�/�"���|&�[������$�� &��֑��+��?z�S�L�|D G��˟�a���
�=��►Pٝ��19����l�_���icU��5uPv�N?G�|���|V$�m���i���gz�-�Pj��c�����V�X>b�/s�2e��z���W�E��C2'W��y���s��Tb�9�?�ݵ�g?I��~~�茉�c����> �`��:�,�Ⱦ�A��0�7�� ���9���?'�	����̎w�����b5X�=H���}+�_;�9?��0"r"Ad�e]���D��fاz�`V�b:7��P`��v[�à2��un>�;V�����۞���!d`|ޏ������N%���A�w��U�#G����� �8A�E~��V�T��>�c�s��u�Ć!V[��������T�b��8j�+��f2M�ś��^�e�.��
���  ���Չ�iy^���k��h̄��D��u7�����0cV>�8�-y�q�C����X�w�Fb�.���CE�KF'c>���W��-qA��Q�X�Y�\��4�,�a�tq� n9%�;p�I4��_��՛ԇ���˽Y�*��Ȝ~6w���P�\ŗ��zȱ/P�אq�<����?���s"�������ΧQt:SI���4K�XqfW�Gb!�����#�-\}hI�?���X�<����k�H���v����6��>�s���Ch���������n��``���An����oJEh�.c�P��SԲ���<�a���J�79v�%�5�j�V�z��A�|.$0�H�,�`�Bb^�'f�>+cU�����uR��!�D{��p���"��н��G�/��j�J?���>\��٪���~o\��5�������l	����sp�	!Z��S���J��d>���z
�Q	��Ϧ�f��Y�ɪ'�m�s�8��u�9�K�<5-_�c������[��¥�������%�eF\L��7���E�o����ŋ;��樎�JG��Z�~V(H#�����1�1�:Q#*L2�=b찧UP�_�m�K�L��ܧ4�^��e�=�b��)��-�P`���gڦ�tbj���^�*�t��=:���p~Sg�?����_�w-����yHr������:�A�X��Q���;c��#HC�;!�]��2i�[��� LHs�Y
�B��ǎ���bUr��a��C	g�8�+CA'IdDڴ���G����1L\kg�!ArI2DaA�h:��{bDӰ��Li:�-�N���%�RO��)4���A0������	����"n뼐�!��K��lg�	Q�%�&s�l�+���QK�x�04������8�a�<o��tD�`X��9�\���= ��kG2de��cF2�H2����LT�t!-%)<��^��+�x8Ym����GL�Uifʟ��#����%����!���HSN��l_���7y^v��ԣy��^�2��}�?�v~:P�#N/�{��i����������X�Y����6�B+t��i�Q<�諦~�nUO|��H����q���Ck�4T�������bi%�z'*]���D��G%�0�9�T��E77#X��E�h��jO=�������\Ų׍�[�3�u?sE��
u���:Oq1���=mO�
�z̹IO�Ջv7���%�:�|��q�@�!B	 ��4�+o�� �9�<�l�PCm�R��^x���_1�O�w��Y�<���!۪��H��ۢ���!��RE4�1
G����T�W��?���һ	%���L&f8е���0|p��Y���!�I
��S�>��G�*CHp)5��ghS���c����ǎ��E�.�eq9�x}�QjF[粿~XĘF�S�Q������o�+�ߴSE�_u��'RZ����bf��&=r������U}W��W܎�Z�(��|B�v\�8ls3��q� v���<5M��3�
����jE��ث�u �} `���eW���Q*��:���ËD!�粰l��i�X����G�����f�4����C���q4+l�PQ��� ��z���(	��{�= � ��@@�>��� Bj����7�»-�d�A�[,1�g�#�;օ�ǽ���V���vbG�.u�Q����4�!ţ��M+��O�9,�Ɋ�����u �� ��S{	��?������+�巓&�^8Nc�g��Y��-r�̧���{����s]�7ݓ���8���ڶf�l]'��D�e/�y9?[t��6���1� �+�8ջn��|�!�F\d�^vx���q�Y�M�y7��A�GUy��l켭C��M�~wɀH�/�;�Lɔc�ĦRc �])C(= �c��D��脤c�C�A�k��
�S��X�ms�yX�dL|��/e9a"ru*J���m��NSEg�R8$��R��	<A0�̳6���B/e��<�1 @͝S�2���Gu�����J/�*fôSc��"�� 5��G��D�nǷ�Tr���wӸg@|�-0/.?d&�y2��GXmVtr�F�8~�N�����Aw��(���/��:���E��xI!��EJA*��ӱ[r(W2����� A�;�Ǔ�����'�ំ%�4�H��)8��K�@;���10�ӟ j.��헍��4�#*�h	��)��bn�/b��v���py�>`�{9�Q�\ib�pF�E�^��c�n��VڏZ�3i���U%L�����۾�'� R��.�^����#�&�&`��h�ݒL�������0
�а�<�ğ4�]���)̩it~Ʃ�)526u'���u�z���7Xjm�ZJʢһ�<qQ�9}H�R�h�w�� ��I&W�� �u/S�8yj�e��m��{c�`�g��A���1yD._E�Qaep9�	�]���sR�B���m�RS����y)�W�;�@�ָ腋G��*�"���9����y	f���e?�e�q�B��!�RCS����~
G�TGƺo!�P_���Q8�!-0�Z��y;~怡��w���pc��B��a1�~���{l�V����0a��n{h��,�2jR���B:��6ngIF� �iU�GeG��
ON?`=-��������o���i�צ�����-�:�܅f?�B&�A���ɯ��FzK���'�?��;��� �h�E�Ra�<��w��l �F3��z�E��!+����h�
���H~���&D���b70P�%� 9�m/�=`&�B��5��{R8m�̩|VN�J�N��(W]%�+cj���{G��f	ׁ�}{�&�R��n=y�D-��5�}���PS��ѡlp]Z(�N*�+�o�[�~�P������	�J��h,�dK�W�.	+64��Xg~�O�Ȕ9�f�\��4q��?�D.1���W�����eVG�%!n��É/5� Qk h���p�����󯬇T���i6�n7L���)�"��%�nl1I�^eg��G�����e���+_D����Yfgq�9��F�,O.��"b��X�*>�w�]*��L�����hA�w*��?���x@zj���H��"o�	sX�?38���!��;:�E��T�c��Tn���&�ܷ��m��I`"x�	ǰ��0瑹LJPk�ӣ�}��+��wx��*����w���LY��k},�:����|色��!���SF����Si��.�A�3ʮ�ƫ�U��s�}�v� �y��?�IǇ!AZ}	��Ea2�����吂Vږ���s]ܥנ��D�� �}�cĪ�\��}�4���ġ�s٣!��rD�VX�1�F/���  %�ǚ���K=5��/i\B���JK����ׁ:�lm�(���R�>BY�N{��� ��:��_	��0�@~�W�.]	�o�f$��u�Px(D=A��Wy�B�t4��l�>+<>����K%�I���K-�i�b���Iɏ�әw�3WD�g����=��ꉜ���J��;�z���r:o(V�`�T]_Ц,�#�q�#2�e�񼘢*��
~��4^VaS��0Ȉ�ܻ���c�U�zhW��!�t���(�{e=L��2}(��ḏ9��lHrl�Od}m�A�F�s.�q7�ǂ��Sc�������6�����Ȧ�N"�t���p��E�5�I�n�y���짎��a	���@_�++�hrJ�ȿ4x[��$t�S,Zx�����67==S[xP��5�I,�gLޞ�}��N����|
�0�"[����]�`9��}Ř�P��$�-�W�8��ſV��X��Ф��=D�ª��gt��<�Oٟ�5q/ ���`�
�U�RR�����ez�x����|�O8󵪾�T�6;m��"�/�m=|P�`��,uNϐJ-FfI%IV�ɊG
܊���h��4�V5Z;eЊ�!,��w�o#��m�J���%O�⿴���f��H�8`ܜ'�%�����ʦ�G���u!���ƍ��Dt*��Ϗ�O�����떢��q	"����Kh�EEt��Y�9��:h*�h����n�+v)���?�	>�@�)����*�y���5V{̙���kXw}⏡����z(��&d<����ɞL�]2��?���HHѽ����D�I��H �}�jB?�_�N�\�W��f� H��7�?����w�3�Z��	�FS�_��T=��a�K*W cv��^�U���ԙ������5�_³vE'��;ف����;:;?++�H�����Ʋ}Ch�ʬ?j����
�6�F��i�k�}(������@J����#�W'w����j��PnK�q���׏i��ys����;T��<)�4�#���e?U�O�E���ҚX���7v�� �R�<r!qEW'�O�"�$��5<�̳,�F1���J>�<��h`s�[m�.������\�A=��?F���Kf��޵_8�������㷌׋ť>*���r2K��vF�6��|6	�+���^ʭ�ߘ܅xg6�dx�x�����Nu/{nw��7�h��g����UC��(�1w���o�kyHiF�x�03�����ud��b`ٓ�S�A��|*ar/��5Um�6N��:�vP[B���}H5��g�8��q�\��������\f4��f��p�s��UXj��8�x�����րl��������VD��N.�$a�I�R�Q�{���W&�����g�����%��WW��c+�D��B�����st?w�H`���`t,g,�[`��i��<�'Ҥqw\�e�
|&�_��)���d��1��4oNN�H>85�R�l��N�q����A8ί�3o	��\�XlȘ��T;\��6�������I�N$C̙��ǐ�3ī�i�7]N�|�F�8�F3ԏ�C��Z����s�t&�����s뽺�<�)����8��m������h+�2X����K9�������+�k�wY�x���M5�'c�4yӡB���A���"�B{D����U�=!6lO�����������b���$��j��翠0�V�� ���`Z(`���$�4{zC٬ }���_@b&��oqě�n�M^-�?Z7]�B{��;�'r�9*��**Gu��}��q�p6�Ґ`sjR!M��n�#<�ɢ#�2�|���%g�5T�WO�bD����|�~�ð�$��v�6�c�a���q�D���Kc2��K~��XM�����&������ G��w�%}pIEu�A5�����>�	\� �'��M�踉�C �6N6�?$b�^j���;����t4,fT�a-�u�HR�U	���O�b1��x�r��%7K�v���Yi��~2fH�]a����t�n�V�]���by9�w�A��P-�f���g�t`s��N<��r@��	g��c:gg?Zuc�/�6�T����~sME�� {�h6ӵL�G�03�ƫe=F�RYޱv�[
���<�E'�6���{��Q5x1��a�l��.1�yev��7�RC�X���M.^d4�������.o�U��2s��XPR���*�0��N~)�=O�hʡ
����RH�yf�W���Jc7�@���#�+���n�C�:�ulX�v��Xy@Qۏx�,矠XX���^�
�&gn�`ZR#B�9$��jP ����&�3��AK��ϝ +>5�ʩJA��ϛ6ɓ�u�ҁ!7+\�JM�5��1�C������֑�h쭾��	��i�9-^� ��cLZ�b�eۅ̾5b!<���2s<F���&Ġ����]&�p�h�|_��Y;/�+����mSp��9L*��<�Nh��σ�hhӽn[s9,t��&w{�HT�����?B(5����L>�Q0��"Ӝ�a^�>fR�I���})~?ܽ�t�*�%Ec�}=n��u�謐��^�<v���7���C���x���||��X�?�8s�=B�I�`��upW�yd#!ǥ�����(��9^�P�8���m?f���.���7�M�ΦZ=�Xث��l�5�ÔCC��Z�!n�]��	�q�`et�&Gc���C��s��J-��A�9�b�~M�H���t};�7YZr����E�_�uC0��6ԲN,�����㮥^�TH���}�S�X\uk@��]<�\�?������bP3_�����/m�JY%Y�_��T-��v}�.�m�s�������z���ֽֿ�����S�L��N�=l�x��-I� ��{b�1�@I������֕�������H0Ӧh,5Yqb��R�&��L�H����N~�&$A��E�Ǒ&o�Ĕ5.����nYv�`��m������\ghf�or�
��bRF��� �:��{�REg��ұ������3C��p���g���p��ك�5]g��ڳ�Ijq�	���^�s9������>M=��Nh���8�Q� ���Q���C���m��&GkCqV:��������u���ݒ�ޘ2�Rtd��?��U����2�DL�dQs@��.�A�>�Ɵ�ݛҺU�Lߎ.g"pjƍ���&�t�	8��	�'�֞�uƧw�N�����ǒT�+�,\�	�2v�ԃ���K.)��f���C����o
a}`�Ta�}6'I!��˝�^X�	�}�N�AM�e׼<�ZK�p̌�j����>;����t��tB��1��N��M=���R,͖{��,�!S�ێ!��o����D���!�����~h�c�?Hc��ϟ���m�_D`������rT$)m�z ��+e^\�-��)��P����y0�`ܮ�%��9DG��.�V�ߨ��`��u ���zIh0�&�na�R3@ �\�0Ҍ�h�����aj�nD}�K��{��Q�3�!�<&�[8vO�b��XV���/W�
�.�SUh*-�o�P3T�Ӗ� V�Lл�'|���Q�;���<�́,�
�9��:-a+>��ߏ.��;���^I,7�P�ƌ݂�ErxXA�_[leX�u��` Q�q�����-�H�s���>y/�By|�4���Q�����c�$答$��B��>���N	X�&�oj3�K�"9�UM�o�)r��Q`Eb�]�+�{���2�:�_�nT��CD6Q���Ǥ�Πh��U��$��(NṆ�X>N�^�\�bKeӈ��o�[�^���L� ��6�F�����>�\���$Ü�$����Z�d2���;[�rt���hz}���x��/���ɕ"��.f�)�n��	7	e�+ח�W�%Ŷ�-F�.��m_��tD��/8�	á�&�b�ξ ���Tj��w"����1ۡv�
�h�O����eM�6�Jk:�o����>��H{�<���a	��_��ߩ��e���������1��=l$�O��K�:�K�Q-�`�^���SZf5��V�Z3>t���s��	q-���s�VH��&)fm�*>0�}�M�pL�_�쥺�h���P�!����,�!�8q<���Q&O,���v%@��8@�[�6eq搠�����s)4��.oMޘR�$��Wn��w�^	��v���r��d�0j�M<��&�H�S����0tM��M����.�X����`@E*�\�Q�,�	�y44'|P�����V������^��__8/���^��:!IX\�5SMPS�s)�х���ٻ�d8m���?{mت�iԽ����礣c��ʅ�{o���;�A�ө�OW�es��ג2p2bQ�<�u���b������9g�,�gy]6'�`! ��{��	�҉�e�ѷ�l��[D~{����Җ�Z>��N���1��n 
��M��ȃ�i"�5iN��Z�V�vG����k*��s攄��B)W�E��'�Ӫ�>��5��6�4d�m)�̍�(��=ɷq�>p�/r{������k�M���L:/o0�*viNgp s0'R�)Zȏ���"�9��+��oݓ_��5����P�@�J����Hn��@lȂ��o�I�p��DHWJ����^��7���W���1I�0��."a���*�7gk+V)�d���k�c>C��y��.����I Z�X��
ş���h"$a�  ������ ��󫾑7���$�j�-�Y�K�B2ld�|���"j[uFxV��l��¬e,��հ'&��<�x˿���!/U�#<P����dm������mH�#/�kl��,d|�y$C/�g���J��7�]d��v�o����@��G�c<��vI�:$Y��药�QUd?ݶ�B(5&oFEVVM��.�H�m�6/#�fF��k�\"|F�'��Nm\\�$����,=�|b�S�e�l{��ӷ.7���b��Õ2���[d{h�ܱ��5Z���̏	<r6��bW�@`���VU���nC;�@z�+nU�������$��Y�0��Y��բ�MغK4JO`����_����������v=׈x>eeJ�ͥ��mg��^�k��x9�k�[B�Չ��m����&nm�&�D�<GF�Î�H&�TO���/��.9��=&nо��sy��`�L����S������A�Y�Ć+�1������!��y}y�sb� ��')}��_�b�Z��N>�A�=(Õ�M�?<�=!r<��aR� �J�p�k���6���>��Ȟ:�!]���!�F1F�R� �.9�ɷg�N_���N%��JDʂw,z���qǜ�#wx���;��L��m���N�o��m����u4E�u�,�V6	5��U�.hȤS0ly��Ó�e称�,_�^����
"�f&��T�D�UĿ'j1E�# ��2�[����ˁ~2�aq>�����z<�4P�G�=~��2*�	�W�<��z~	q*��y�Ɯr��c������~=�2���S�3���?�Z����|��O����)��#@��h��C5���i /���j ҙZMb�nc�E���v�^��=�R�t�� $��S(�,4�i��e�����o�~R2f!iy�����1��!��T�(c�T�j�H��w�^W31��Au�+�_���Yk��[䘘D����g4��Y-".}�.�U�fr�-��q�@~:�)t�U7���A�%$7�!r|����Ym��ٴ�z2�4�;B�,�>��p�moMHg�u
��^�y��On���L����U_!�4ˎ���A�d�0���kB�?i���!�h��u�]��QNM�!^��`��k5@�%Lk�g�!S%��e�_���B��᫔�52T����}�ǳ�D�e",�D=�4���`r�q�~C�5��[8�ļ5�X�{��	�J1	���;��OJ폟��D5in��M�}�����eu�����%"�6���L-�)���+���K��,�@����LrA�%9��~(p�j�S�0G}��Y�o}���DxO��MN0�[� L�@1��%�.9� �م�'v�����A>�*_r��S澍U�;k]�����P�җ���R|H{��R�l	z�2�ߵ��q	[*�VƊh�h/�e���,D�Jë�e�y\����<;ᎀ�&8�7���#KV}F��F����IRzzd�	���I��2�GJ��I��&>Q'��j�4Y.mw@�����E��҄�PxF6��o��r�1>q2ku��{��z^�4[m��UA�P�[g�g.��?�R|���J���:HB����_�����`����%��Esm��5t�<��<���3>O��%w�Ն�]�v��J{��D�L�RVE�>��`O�N�d��}�e�QI\:�xYm�b�0��O3.����c��-K�2e`E�|TJ��c�>m�)��F��	���*,�A���b2~b�l�|YsM���6��ݛ'�wP�,�yu�12�����0^��r�n(Xr��h��	��9�~0��0{YkW2�I���H�6/���	�e~��V���Y����5��Ns��5�??d�~k��M9-l����)�+J�T-�}�n���*%?���S	��B��� �4Y���H�eq�t�����٣s��W��Z_���M�7��UW���w+IEf��U�>����BM,�f��s6��`��~��Ȋ����I����!%�[t���e@5g2K)�2���K`E���(z-��:.�,��2��yQ@	��?���Q��r���j�P��(q=6g��@J� �j���ޝz�w*p�p�1�}�j.�X�6��٧�@M�3�g��a%C��0��ݘ9�����B���+�k���������QD�t����K�.�z)f5�N!�Bk`Ўj�w��*�Cy�:���<��F�9ׂϕ!u�l�#le7G����P�������w��(MY���|	��ru�GYRx�.Z*�)�3��r��}&�6�L�-�
A����F����������3b"�JΩn7a�E�#��-�|�ׄأ��*M�1x�=ꦗ�l���NaTG_�U�p�K�2?�_��$$��R�倁n��=�j��.�q�t z�SZvA}r6�}C�*���w7��w�sG�l!�$���$����>V�o���w�8��4m��Bz:�kʍN��r�p+�Y�p�G^w��@��p8	.Ηx<��g����o{)���jvK���U���q�s��B�9W�;��(��o;��I�N��Q�b�%fM���+��Y�<;�6x;��/�j��[�	��Ԅ��D����T�qq<if�A�f_���t�]b֌�M�\�5^e������B.���A3D����7u	����� ��F��T
kn�cEG�t�1�+��:�����ڮ���;��!�d$��N j���I�Lpx%����a+[�^%��j=E\θG��}-�\3�f�,�@�A��>��^�ŋb:i��5����Ё ƭ�j�-j���OI�X�?�p�:��2�i�
M-���1������zF#m<*׶0��
�6��
{э�<�0�Jz�F���u`�zxM_8a_�X0����YU%�M���y�����H�聭�j����;�A�9��`�����9�2��ho�`��3�r1G/H�+@�4����f|1�:i����_�8��W �ȯO�~�6
f�Ԇ�Yl��.���M'�r�_T���X5�f�&����=�O���+��(����:r;y�G��gy�2[d�p�H���\��L��KUe�,�B��|�(a䣔��'��ɜ>)Ud���|7\�5L�_�� ??N�4o<�q���Ye>��̬���,1�j!���hG1��J��F��L���6Eb�.�w#ǝ��S @�V)�?���I���D�˙����_,����m��-�~�D�G0���M��٥��a����S<ZF+��������8߷�}6^o��c�yD���4S5J{'޺r�P^�w{}x�k�)��Iڠ���#ǯ����)&Ĝ?]J1@�=�*��#�j�m _��v�S��G��� E�����n%�n|6;v�H���	��Y�1t=���Z@���[0YB��c+�ま+	���ya7���G(�$Hc�� ���І��Y�!,̳������Y�_ZB���yY8Ŵу�B�mA3����_R��]c�#S��ܱms��*E��D9py ᡒ�*��IͳC�����K�%�sݻ�G��mh ٢��v=��"/{0m��4-��].��a-2�6��R�)�W�Uj�ݖ&
�L�,�d�U�Hy~�TW�]��߻4gp�T�C�ʈ��>��w3H_6k�yH�w��=�A4!R)�A$YTPKO8\u����~��b��Z^)�a{��I�X�y\t�Cz|�D<]��{�����[W�Fut���3��~�~��8�����ˉ[{w�����S&��wUĶ~���p8������_�e0� ���/�Tͱ���hW���x���\�)~ �k�[����e���G��+����N����}���&�9�Wc��#0�� b�q��v�6�hA/u���B	^�6SA��D{e�|�O���t�rQ�$�%*����L�qteL�Mܟ4z��+��Z�m�G�����΄CV��0�Is�+6vSp���É�~�Z��J+�9]�h�DP�آ�+���_5)<�Fq9�V�i����}t��P�*�1�^j��K�t�QC�$���ɓ#x�pĽiR�jnnB�� 2H�[�=��:Bۇ{[[�S6�m���P��E��͖�L�M)j��`_� �z��������ZW�v�wu�l�Jb? o�P�n؜� W��5Gg���j%�P==!p���K�{�a�, �2���ŀ�G�o��`�i���X�s�?���c�r�?0q�]}�9I�xT}V�Ƕ��.����=>���_�"�B����Av?.T^��՝������
���6<�G�e�w���:�B9]�#���H���������j������/$ � w:�U��C���Dܪ���z��pR�/=7��Q� �Z3������8���&��ն��	.V)�R�J�6��3�g�LPBqT���	8d7	ӍQ���|~&����U8�z�Q�XѤ�ԛ�V��{O�pO�x�uu7 ��f������l=��+ 5-��v��&�Xd�=����U�~�46�S��ʑ�ݴ���6{��@W!�3>����̂	�l�]��ұ$o	�n�0+�t��DQ�R����n-֛���?x���[�d4�LM��������e[v���&hlF!(��L �/s��i� �:����׻<�����6.��AB9�VR!�7�&ܰN�v��2���w�,gj�x�[�������S�.F���%��O�s�����_f�L�2�m������|��a_ʄ�횿n������œ��,7��|)h6zy�h����C��̜&� \J�fV�s���]�be �}"��i ��/�v4�$�t����� (U�(zB1����c�gZ052�)ӈj�w���m18_��A
$u^`w1��o�qX��^φV?��<=��1�*�a��8�_��g��F<�KW .���̖
3g��BtJ�MB�	���@����>'��* -y���ޓ�^�d1{.�/N���O�t���1CC�&����}	����1�݈��21����b�哊oar�O������-��3g��v���7B��a�|/pp�{j�� {6l�Ep'�@~�G1��#��(�n3P��2Üs�~e)%d�O�1b�!Qg5dg�\�Le�X�D��t3��zk���*y1��kՄ~j�;^�9I�IR���F�(-o�F���,��"^�s���8��
մ�i�o^�Oi��PV�d5���u��� �j���)�5�t����	N��Or��)~d
��^m�N1�C��� �j9rZ�ې[C_}gM,���^W(ݛ�@�� �45t��N�<|?��|꼄�Q��c}�����p�hm��C�཰��#��+Q!�o:e�L� x�>Q�:
���&�b�1�jz�8����t{l�A/�d̃O�oB>�Z+A��3���W9,�R"�x�� �Lh��ڟ"Ԃ �5�{��U�
�lA�`;}�=B2�3���R��Ig^�b<^�Ĭ���e?��!�U6웓�M>�.��T�\i�n;��C��Pt�ܜ����'>���yy���S#G4fO�g|����6�}�\Ϻ.��|�:�s��r�kyu͂`CK{d��v�1Np�7��]���4a>?��^pہ�h�5Q'H��4Ѭk�N���G�p���I�d�W�R���G���V��������U�>7��5����_���8�ᑬ�"&m?~a�A����Д����~.���U�DSrSC6�i?�e��"�Ǚ?o�b-�lg�`���&B ���%ʒ2Ό �뢽����"�4C:���W�h^4qZL�f]x��L�z�K;��[�朩G�d�O�3�Y�b�����:��H����WYgf!�iVsL�C�>���S0�D�cԪ���ځ�>�p��r=�#����C+���v�Y�O�Ol��p�G����6��[7ҕ��ދ�/��e��2�S�Ɨ0ګP����wJ\�z���E�s`�=9-%1��S�����p����M.�.��bq�f<1u�����틱�,U�p���H�oDB��h�����l�ዣ��W^��v@!�ȉ���d�)��ϐ>���ٽ�51	�Ma�X�I������&9��<�㌢Dʽ���x �E�{�J�G�`�]3X����*��;?��NI�,�n�̓ƥ���_U�t|�����HcG�4eA�u�M��/�]���{����k����e��S��5�@j�rwV���b�h�n��#��{�G+���0K�y���_�C_���_мr����hB��{�1$f�p�� �C;ȭ{�"����g��z|,,%�FR���U�Z����Ʌ�+��V�Ұ���gN�m���|�E�P�������q���Rs	af�M��Y���;�z��l��7�rϓhw/�����F�B�$D����DEO4^s/H�!N6�۸�2��1����Et�;�� ����ͨ[�pp�γE	2s���{�+��7���� ϒx4XA
��i-���u:�Ah3�{���@� ����Ϣ="Sa�y�Z�n�n��Yv��vi��J�Q��	ni�}��"�6L�ܟ������ه��G��&�Jy]23�FxX��ݢ�O� �`_$�u93�ψ�#}?���`4�d*R>��_S;"u�͇�|Q,F��Y�
��2;�c~��n[}���<��d�殢����\{�. �3��&��õ�Q����|�nAI��u�t;e2k�a�Gj+�E);��a� "�.�t �4�ly}3��I�c�nQ��LN�>�QR�ў�S�i����H�t��v���:j���E?d�8�ԭԂt��҅�Ӕ� 5d$C�Oͼ�~܏�FCW��r�y�V�oW_j2~��*�� Z�7�%��cp-���sN�9�]�a������sA%��#��#���Stv���	����քy�bS"�˓�jZ�9ϩ,}�����}�`.�o�uS!��big�m��Ԥ���O��m��	KNG��h�-�M�� &��9[iB;5��hsk��;`xǁ������èP����Cqu�;��n�:���͝���`75�|��d^��i�F�?L�x�Ľ�HŻ�S����S/V1Z��+.��OP����ҵ���5�o8B��q7���%Ȋ�v��QJ�g5Wpc�Q;�\ﳤ�㬿�h��hXz69AWYc���QP������Yƪʧ���9�T�w�!��y�H�?��t�D_�2���	��S�P!w^�S^�gl�S�CqE��P[v����:���R��{�ZR��Ǭ	FV���`S���fz��6D����^̔�'[�%s@�F~5=����c
��|-/���Z��l��돐.�f�0�2��!�BD/�8Za��\����j��n��+��	Kq�5����H������*m�{�����>X�!Z�~N[�V+��� �6#��?wL��E2��`K�aG�qs@Uc'���	��pv�jym]e@<�&�If"Ml��wa���p�H��yN�u�wk|/�NZ%Nv6��l��ݖ�fߖ�t�T��J���0d���P�-e�����d�YO��4�1R��]
]:�T�N��I9��$���c���!���EW�~f��r��رAMT�i�P�3��݂�q�5Ub�Z{K_��J��aC�[�z��c�J�(ޛd����2�lJ��©[��L*�M������i$I����A��#	<�]�:��u��]yw�s%*�� !��1Λ��Z��̩ �% 7�R��Pw��8�+K8�<d>2}��a��+J��(
K�q��n�I��6:�v�Ӝ`��Κp:ύZ���.���`�- �<��U����,� ��E�f��:��1�U<��̌�Y9��b.;���b�r��԰h��W��s�5�D|;�%B�>�}�*Z�EC��%�����48�ZHo�e`�I	�{����z��*�M�O�z_��&߅��`Aa�*+:n���r���xa/�D���ʎ������8s����B���:�M�Υ'����2..��y���¥3h�A�_���r�Y� aB��A����
��n���ش;��#�L��a��hG� 7�dG��8T�o�/2���-��\Y��V9��P���J|L��}�*�7缲�ܷ��6����D�{R�G��P����aPO��=v%����uj��[G�V���-$sa���J�\;0��%̙'q4� �gl��	�t��������=��j:2����
_1_?z�!���=���H*i��}yo��f޲X�Y�?���H�USkJڙK����}$�� �&�ەj��U��ν{�f��w��{!9#@?f;-KA@=╺!���N�kѓ�\��&~���ރ�ʟ��C�E[��+r���e)���su�,
�g�ߓ3Y��g�X]��7�2V�=ʦ>�P��NJa�Mg|<Ő�o���b��j F��2*K�{�#P����?}1�3�5�lR�KXzM^>$.�p猌誙�S�c��S�O�{M�S���}U�অ)իR�S�N��j+C �D4�@\Tp�(~���{���=���\F����F.�����j.�ڗ�]�\�Á���_n��2�0*]�:[YJ=c���#��Mo��3���g������ܚ�%��`}��G�{:����J��ŬX���\D���y4�[��s����$NM�/���dK�������xiQSt�ǹ�a4��(Њc^�>#d��O�-ɤ�6�X|t�<ohC�ٜ|u)R�	�-\���@������s�ÎZ�"I98M�FM�J؏D����j��Q���3��X�40�6�xL=x���
�>~�M�J�2�y��<�BM� ~+6����&²����ܿA�	�YL��)����,T����a�'\stu���ms����ak�7��I=U�'�����ˋ�?#O+�fC�ҵ_�"ms�Ӯ<��� ���!��o}�����su�Qv�x�<2<��D@�Bm�n-�F�a�;yz����9�[��y\5��A|+BM�w�/��㿐-,z+wA�_�P���K;���� ��V �ݮuc���H��'�%}Ή�C�%.%Z6�:�-��1x���R�<!p���S��^�0M�Q�EqA��Ԉ{wͿ2D��r�>���u��ޙ��H�U�%�k���(v��)��'�l�<��:�W���3�����;��o�D�Z# ¤�2�Y�{~���=.¢
���Kl��\�Ƈa��p*��pk�K�-P�]�x��ע�T؎8���J�"/0tv��]��b��i�dO����h���E�`��Rutbi4�#�ݗ��{�z�O�1w/��7^��~Ӳ"��Jg|,������F��{���@sPV0v.�Q���g�v��;u��E�t&�p����=\�0�#����r��z ���cbp7�F;)/m7���j\�/�����E�<|qS&�Yr}W_Ւ��Y�[՗/��RK�~1�^̥����<�JTJ��l�K��G)yq`U���on�X��椢�B���W��""�bu�I��K�k��T�WK�VQ�"2S�]R�9æ?EW���te�y�����E�
�g	[�K�� juK�"� �Q��M���Ӥؾ��ٕ~��@���yU/.}$ɨ�0a��㐻��Gك��Z�3����2,^�p���!�Zw�o�6)xa�L�xX�����1��T��*����*
�^$�?3mH�I�|��R�S.�K�Us��� ��9w��\U�:�:/�>fe�\�{4����O[��G+�ҝ�� �N ��2T�ڡ�v�$x�8O'���{CҶ��p �a2�؀Yj8NZK�ڌ��s��Q�|L��&:;�f�r���f{4N)} ���&�P�'��
N����>5>Bo�٪��e�[I�ڏ?B�j��o5sêkԏ��ԧh�5��3CE�㓘�(!�e��t�J�%���NElG��n ��{x�F�Y�ӁUux���Š�;���ߩ��fy����<�Z� m�L2���)�i�ށ0	1�
;��>���aЁye,�Y��s8�S[D[w�u��ݵ��yS�O�Sl�Ħ�$����Þ���7xV��J!���]��c�n�����U�b�v	<k��J��M�5(��uu�<P2��67�It�u�s�2v�N��0U���v���9/C'Ze���:튱���]o���U5�?93A�%ϛ�ΞO6���2�^Uxj?�a1à�ݣ���J���5�MaF�
(��隞�4��4��=�J���L���*���������tۇ������B7�+�D�Ւsi��6��@C$��s�|��_3
��` 3���]8ՙ��Q���B����%�^(L����p��q`3�����Cݝz��+|1���&ZK��6�j��޽�T�|Ў����� {�h'e6Q�ɵ����6�c_�B|������|�V��6(��Qjl�����<**[�7&�t� bㅤz���7~�c�����H�cF�e��$ɋ蝟��"�&n��'_�#�P�P��T*9]Kh�w8�E��,�.�Pm��P�qkb�Ȧ�I�8�}�?W�U��a�7X2��kC��"\B&J�����E�\�v6\&�X\4(�k	@��ӄY�ܢ�x���Cw#��TC9�9�6���3$�;fX��ܳ\|�X���_��"u{�b	�������ȉ����ғ��ӈq�8��o���':�U|���ի.�td-謰���\�a�>(��E�8�Zh��o�&�ޟu��a��R���r�49<���jV?��/Cj8���[ pF~+v��v_�0��w&����i�ߥ���J�Q����?w��1G�`��u�݋#�_��p<Iݧ��C�U��s$���Usc@�`�+6��h�2Sg*1^�sd]�U��L@���V	��2C�O��Sr��T"�X���#������.f���4EhnX%qd⤼��/����M�A�d- B�&���E���ڀ7���dC� �BX=;����;M�V|�G&���L�Q��
��Ic�IS�VCY*�b{Hi�������ɺp��Z�����{6u �Lw��V��f �f@���~�.I��|�w��A��>'���%v	h{.q��\?��ŭ;Ȁz���tX\�B ]1�8z/���q�Iu�4^<���H���t��j�ݼ�Z��h��Hy�x'%� ����A4�-[WE�URW��H��O܉v��#�N�SHĀ�J�����v�fi�|�d�nQ��fI�>��W#
'���^���,W']ō��mT��Pg��������X�J��x͘#�\(r﫾g߱�B3�f��-{�M�@;�Hh��RϜ�O��L]L-Nl2�Z{���n��1�@X�q�P��$h���,�L�N�	v����d&I0�A2��	��|\��+��1Sxϸ�;���m�a��Ƃ�}M}ǎv�V��������o`��W������ap��W�@�f���,�A`-����'�/-��L�#+'��y!���r�Ӑ���G��J�f��2�$3h�]��t��"����Z釨�U���Y��Ij�mZ�y�����H�Y����(t�#>5ɬ�m����g�:q��c &��3�Ϭ�n]n^��7l�>�0���8��tj5k29�瓪�1Q��9�`�=T���O�6�tV�#ơ��*���48Á u����4j�vx&�dLκ*��O9��B�o��G�u�n���K���iv^r��5k��(K�h�]U��ݣB/q{7=���[� ��Ο ,�cꡧ��I�޴����bQ?�ݵ���~�IkFe�'}��6����e0ě�EDdR<Z�ݦ<D�*��Ԃ��J���smq����oWiR�pG��oe���p�6\6��n���/*R�A��V�Ue%i��p�- ���/���,����N,�ĸ��|w���q�^��!p�i��]���U鄆�#��S��jo�|��8�YI�A��Y�C~�d����{�7;�+��碀�JbS���.��F[IG�����S3�r��U؋E<�	̼WH�ds,��1��1��,��f˺��߲8���^k�3��d!����s�v͖{����8rQd��@�h͢�SXB�%���W1DK<��'������nr�9�ϣ?��,ޯ�V��Q��nJO����]�
��1sx�΀%�=�g��%�/q�gs?�r�5%2�t!4��rօg�@����i�l�J���/�G�����̘�ƴ��H�xb�%JJ�1���0����h,��ͱ�}j%��3U�r�m0�<�'D�um��Fh/x�zA���������DF��H�K�D��W������PE�E���c8�1��w�A��B�c,����s���n��
�5q<V6q�3���VX�9�V������F:�<)?�J��Ԅܱ��.��M��y2����<���r��ƌ����/���_�**���r콚��G�/#v���q�h�����?�cI�ؾV1j Ο�8ҵ�z���EY6����`J'�<� ח���6����o���GL"����>���|�s��'��� >�\�(�#����������f[��.�[��m�#h�HkC�)$G�I��bD)�Sp�$�C{�n�sn����I� xf�m��]v*UaK�u�	-��H�`r�v�|F�#�'�mhK�#@M��_Qp�7Ǧ�Wd�Ja�B��ޟ&*���x@��<9�=!4�*��X{��o�݀�5A�������-��M/�����k���'x���(-7˽}��0�sxQ���]���Kz������=����1��j�#���(�ڎ�����FK�_%�v*aԚ�Y���^�{?cG��S�]�9��Ye #��e	ޝ�}y��H�a{?��9ʪ}'���OL��g֝[u�
z������g�@��C]�!8����� O�c���{�B����3BN��:(UL~҈�͜]��5\����AW(����A���<��Xt?����%z<��}_0~�3�l�l�Q�����q̑��u���s�a��LwP�"֘�������mT�aq5�X&�x�rg9��竀��q��6.V�y����'�P���ʉ�3�ޣ�f(��)~*c@�+�=�&�_4����ӟ��l��p��HZD/ J�_Ȭ�oԝ���+x'�|���>��qK��'� #Z4����N�n^p>Oe�j�l�Ѱ��RaHD����S�0h�0�Q�$΀ Bʀ�ØV�2�"�#�Qt�{GkVc`��~kPe��R͹�P���V��Ӊ^�.G��֑��g�B�����F���P
��Bg��q��5�4��Erq��wF��M��0�A�_U%��lQV�.)yFԶ�����]'��ާ�@c�-{@���*R}�hZ�s=�g�1�6}6`��H"H�Kb�f I���:�&�7����Ee��ofH�ON�y��l�6(Nؓza��J�ڭj�k����疐��pJ#�pw���N�����ӑ8�$pWx�ham��B���ڧƮY>f ��������� ��k
��\W�[l"����ZW�:g�{�F8C������Sǎ�d���8���,J�&j�\jϕѵH��>U�<�a��~��A�Kv���*ùx3+s�	��p�\ F�8t}Β3��?�F�d:~kz6hXx�Md�-
}���#�p���uc��.P��jMNZ�ԈN���a�V_-�B� ��a�T|�������[�'�i?a{��G9�|�
�A�Lm�����s��v���g	`�~9���܎��e�,A�^N�޻Itݚ�Q7���0���g��t�a=e������F��[$V�l�,̌������v�Q���, 3�x�0Bl�m��䨰!�)��IFq���U��8�'�T�t�Y8����!ǔ���H)�iV���p%�;�k͋yK3���������[0T�<�N�n�q��4���]�@8{�n���r�������|�r��3�gV��J8$�� D���to�i<|�K��Ns��F�~5�r^��vׅyE�E�������j,���&�8o�Z����I�W?x��	�5��e��A���{�"l��V[�.��8�lX��0ܐ��媾�����S�ؕgp�;u9hAF3�����2�`G���|��؟^����`k�EGe�Ig$���S2a5����ې�
�U��s2�C��+�� &��V-&c��R���m�|��l��h Ab@a��^+�R�GM�cY)Ze��ԫ"��o��Fg�:�[ �cj��`ϸ��7O�c��8�|���3��Nל��_�v��#Y�@,Bd?k�;�..���5�u���!'����~�P�I3 @w/�th� o��7�&@]�����S��D��	P+�\:�1�] z��(�fD�6��"
��������@�m�Cl��E��r|AsM�ά�6L��wZL�7$�W�|����w��b�>ު��b.�'�=���G�fU1jl���Җ�O'�4�ꓧ�9��3|����}�T=B���K`Iq�'3�����!oz���Ϡ��ȥ��0/P�tN��8!0�W<x�� 'yV��0�ӭ��KX�I�U[!���G�&_�����|癠����9�qቋ�ڕs3�s��%"�Z1��[)Ο�d���.nQ�)��$J�c�˴0꓁y�ׁ7�"��2�s���إ(�i�9ʳ5&�{gC�:�)o*�Xr9��0�ܱ�KO�F	��{��"Sڻ������6'�~t�����kA��J�W=cYq?�����A�n��SUx��o�8�Oz���},��S�eF��L�$��Z#�Ǔ�e*j*h�T\$zǑi��5ޓY�7f�� =5����h�<��*"*t������d��N��:���7�ͫ��I�G++͂������Rm`��@�\��n�%&�勺T���V(@��q�K��N�GQ�GRͰ�8�F��Z��7�צ~{3ß���!�7�ǿ۲K���r�"<���ޗ�d��Ѝ(Q\t>�2�b��!��C��T o�izx	7�~J9?s��~8ls��*�;`Bfٱ��L[� ���,͑+���_�EB�{SGJ��LZ}Kp�'H���������Z^ӳi@�w�[`�W;(�p�\>XWӽ��V7�L���,{��-����F�Y~F^4&0�E�Q0�R�"sHl�3FY����B�൧^Y\����E�F!�������`���j	n�������C�5��9�TQ��&�|9G����.ik/��|����T��b�=	�n%�m��sH�@u�G�ЮB[�T�����������5<�3����G$!�Z�d.��� 4�3������2�ظp7�e��7�B )�2FJ}�X�YmR��iіZ��L��~���R�A���B��������8��'/����!bV�X&i��n#O;��ώX���l�KQ=�yzb=6���X)�N[�\m���)�_��e����/&��@����ċ�A��}'Y�|8b#���#by�sp=]��;e���G�]��Rw	ߝ`�k�����1�N�����"�|�?P��=�s"�!���P;y��02:n�R��7�ZҸ:1��Hth�ə���ic��:C%��'�C�У�s��Ջ v+���ԩ�C�J{-�g�E����T����cl�f��?g�h�<����@�cL+�r��D��
~��נd�מ��r:��7ɢ��yz@²v��.��²,/^� _>�y �<�ƈ�T�R\F?�3ɐX��A�N���y��mU\����?C�:W5t� .���
�Ju.?f��U:v�̕���z^�nmI������=��{=�g�{�>����Lw�ݽ���� �xde�V���ݕ�3����x���i䠇�3+6c:�QvUu��C7ґ̂;���_�i�j@�3�1�p�om�%��W�`�]�&������z��<	��������p���~-"N]���%��G�۞�}����٬}����pm>bW�p��c�g���oο[OU�fi҉�E��)bR$}vG����v��D2_'��&�A�����Ɏ�RA�
�1�om7�B~`&i�ʥ�:Ԭ�M�$�+a�h]�4��%s*\��e2$�LjM�	���m��I�]�K���d)���._�~�]��6%.<P�"�n�b�ߠEl�����7}��w;q6\q�_��n�<n��Ztx���Ο�
�_���:)���anՔ~�����c��^�ϯJ�����`@��!��y��%D��Vp#?Lj�6y��>1��r������������8�[5g��.*#6Y6W�+й�����(c�J�[7���wĦ!\)�����K1�.ؕ�)�n���(��p�Y���!��_�����a�HtM��\*�����ؙ��t�Ȓ��x���1S�b��^1s��$�!O)���W��]��D��O��q.J�� �%�(�<Y��̹�5~q��\�Ľ��({ȁ��Ѭ'n�f����XE$����3�������g�E�Җ|���~Ȃص`���^j$T?���>#�ê��&�M�Ȥ�Si�
�)SR��`���W4������Zr*F��a���NEz:��s�C@1�L�E3o��=R�bk�ݪ��?F�[\I�Ϋ���N�L���-�mj�3����bO�(�1)��,�ԇ*Ӷ}g�zH��8@ؓQ灺��,��t���`hj�qr�Ú��U���6���a��b�>����C�#N����1�����ɵ�5�0�<�пwa��N5K��{:�fo�1�J^GIh�W�]bT�eG��D����3��?,2��.����%�ދ��fF��Za�Q��_�e8�%βg�����o���,<�T�ݱ-��<���e��o ?h�����-��vq�Aė�^F�>s�/מ��	�a���& ������%����ƨ�Ù�!�h]���%���	�H't�w?�#����s��*��G\�l����z��b1��w؊�6ROH���+����J�FQ
{f�un�ύ=u�g����)�j��&@�<�S��C�U���
S�,Ӵ��p;����M�Ettо7���=?��ڨ��p���~���
l�Q��Z}�Cu��T���!2%��Ak��9��ҝ@���S��g)��c�s�#y���}��(kBwn�q��dw���sQX��hX��w��JV����uxP0�	-�	��]���5�}m�,��L<˒��^�U����!��p��揤/���D�x�"_
s�Ӛ {�����L�e��X
O�h��xn��*�����+��/�HN�3yIu�ط'u]&�e�G��klÿZ]=X#aϑST��1.t6"֓`�%O�a4Άd9Ir$e"o��)��C�7����R�&=.OlO���Դ�
@�G���@r�-��0'{eZ���8�l�5]����(����A	+Ȋ���2.M"��"V(D�3*�XW��*��;�˯�-�.2}��s�Z/����Q�<�&�I�[�E�}
�ٮ3.�o��	g���Ѩ_ˬ�L|�!�@�]��m�\	i�K��+�[^!�f$��/�e��#_����:�E�
j�̶6f�G�雮�w��P�uW~MO)t�EU ���a����%Ad�
d�ݦ,@C`Һ $[ī�����:;(|�i�@9�QյI��ꘌa����e�1��V�cNM.�`��}.�s(|�r�����,uMk�I�P ��F�#0#E���3ie��Ž8�G\�CP�<��Ԝp�3qT�p�W�'�PM,x�L����t2��&G,�p�{��T{���QChS0�߽�zT�+�:�����N���n����K�F\_���CE�G�J�zf�'|ޤưo����D>#+�줙�5(�JJ�]�2���x ��b�@/��,�2tstS	ց�G���+5��4_�������в���B�ƌ�P��5����F�u�ֱYJ�ܒ"��y�q"p(�+�Dz�hq�kd����eS)�1
�3���e�����(�:�<I��j泤
�5�����t@8,-hnb�.乤@�'q���a��u��(#��q���?{��֌��՝�J�4|smU\�r�>H�b�$c3e���2�fl��ߒ4������ϚmLq���I�b��}
�+w{��N4}V�
$AO� n%^��+16)[N���rs�xG�r�g�s��gf��|�d±kjT�����ǔ�r����qז(��u�\V�bb��*�����~]R�+G������h��}����]�%�Zu��'�O!��'�\��6���-�D��S=3d��#C�c��!�7Y;m�K�2��d�Q�耛���42;r`m��7{�rb�
^�H�~�G��k�l.��ɥ^'��N���
'�g0^{m��w�2�5�m��1ÜS'@�w���?�	.¯&(0-"��f���KD(ҧi�/��̶���/����!�%w05�N��C�9~�X�b:*mG����m ��zA�?s4����+��f�x%D�&D�ߑ^"�T8������a��k��js�g_
�W���%�QE#iZ��ѹ�	�����l�b*���m�У��<�^+�r�}9��w��g9�@�I��b��e�՘�*W��О���F!�!���&YȦ�R�	v�Z��g��r7�2�Ի��s�D�0��	��b�,��"k����W��. ������&lx*��S��)�k�3�����;e�/)����e�#��?�Ϻ��C<��S?�,�M���I��eH-K�Z�͚�I������rXR��ٳ��w�n����s8��'�(�%)أ�����U9,q�11���!r <��75���b���a�TfQ�ƍ�O����*!Q�:�W�]z�\�EY�.�6%�ׇ�4�M(b��2XGHO� c��5�	wN�5X��B�*9�;t̇JJ����L�3Z6(�� ��p�����*�k�h�ˮ�w�����s��;�v�p�'�:W�4�J�m�F�1HU+Uq?�5A�~�DG�I�Z[/����ڇ�xx���<#�ѓ�[�c!N�	����Ɗ�x�����E�lK*Ypm,T�O�mF���4&o؇�"�	%�k�I&�w�1 a�j����e�Zwr�y{/��p�r�,S�+�"�5���l2�ǟ� ``��3\!�1b�[��k[��w�B�&� ��Z�(_�&��K���/�
�./��#��	�aeAķmV%8"�=I`S���`d�~}[�ũ�3�?t����q�ȱ<�Z�D��:j�A���0A�C(z�W�s�qcj����NC7�ed�pG;�7?]�4�8�KlNo�-6@������Z�LQ}�|�o�Y�HF�t���2 #���ʢ���r��J1m$����{�τr�v�0��)�o��Ɔ6I�h�Q�'UBo�!~*��@W;E��7��'�Ar�e�q��_��U٘M��zRqӺ7$h�y*�~;r��E*zW�z{fw��V@�y�9�VJ�Ba�&x�����0��A��9��Ɂ�82��,�~�������"��i�ʪ2�4��F���̠:�ܩ0K�`����DÃz1��s����5]�9,�@�d���y{�$�L�����iԡq��_ҡ?�6�)8,y��~(�Wr�����ɏ�D�a"~��/��MX&��kBc���W���!���Ob��9���'2��<BM�.���?�{R5���Ӽ���no�Y�;�*��}CJ	ɬd���s�*��&־�k5�������RO|_�T0��oݥ�<��{�<��)9�r�\P��5EM�H��ZA��x���ҙ�u��QF^JN�(��ո�F��G�m3V�hyN��[�*|���!ŻT�{U�.���:�-9���>5�͑�����`���[���h���o�tkXpĎ�\3R~��P
l�lV���;�8��b��̛���FlĄG���i������{r�7ŧ��F�_����+�JA�݅4�Y��qL��qW��'+�z�A#�_��g8i���ǳc#H�Ƀmg����%���w�����1��'L���N��O��h1k}���g��w�FFİh��zPVP��4��qY�����7�9W�}��/�&�ލ"^�D10�s��.'n. �	#p创Щ����݇$qy�|7�<p?�f�>;w�~������V�<C�#k#;۴��a�����S'v��g�zOVK+C3а8����!��!�d�_^���	!"�Tu[ڌ�
���k7��h9��{p��w�4�9�{1�����zwh�������F�K�x������W'֥�}U� �����h]�l[X�2�7�g^��T��_#�O*��πP�:f�p���j���Lp>EvE��n���;t��HY��t�v*�<����w�߫h�I��^Т~���mQ���� c�\���NO�6��.Il�Zi�r��w��{x��+2�n�`�TS�R��ҦJ+jp"���'��%�8�3��4
�Lp��@l���ITI�|�į'Ҭ�{���	51�������9Sh'�t���rP9��m9��G#-�/�mJ�349��Ѕ$G�/���k�U{ɗ_���`zuj�٧�Z���TKZ_�y�w�dH����z&!������f�]V�����C�A�̓	�Sf������O��ꨡ�=��PĂKT[mb\\��hJ��M#\x�I���r}0�&`��hh(��?M���b-����h� Iϳ��N�E�By���K��.@���Q!!,)�!0OG;���I�f�#���[���e�ʼWϝӅq��KpH��%�.�S�+�cG�����%���,j�C�F ���('��xS�V�>w����" b�	>	��՗U~��Ƴ����h���^Ϟ7Y��2�ҍ{C|	�J�:$L>�=b�LU�D�o�-8{@��ޒr�?�C �n�3��6�8~/[�LLD��e�ՌAӎ�{̒�Yj���<��c	L�?|UJR#n���>���0V�-,9Q��z{�?l��&��L3K���U�YOO[>��#���F%�5�JW5�|j�]ص��U�fN���?�D� /������7�(BC)��ak�C1�=g0%�Cֈ� e�-:�;`�*l�	�O�M�se�c�ТYL8Ǝ�|����K;!��bX-�S�M 3���Wv����'�p�yc%@8�O�[�(�^���s�xK�RR�: ��׸B�X�2�@c+��ןo4��_���@�ސ	�����枴��0�"�@.���a�v��F}n�aN��i��1���5��E��t|]�3h���4���~���n��_h��6�j�X��F�=E����h�,!���I#j:� W���0�O��T�q�=�X�;��DhC&�,�� ����Ea���X�'�/
ۓF&�b-�����6���N:o�(����ϟ>>�g]nmg���=�?���ʎ��:�
�2ܶ��7�0����>�bv�p,���RMF_���]3��۾��BJu�Hj!������+J^9��F�� ?���؂��}����ҤY�Q���$\�C�>���
�O�}�(��C7�|�ͬ�h�>Ĩ�D�=���i�F�̞	���0�b� e�F�S����d�2e�loڪ �� W��A缍[U���ul�h~?
�*��_�X�o��B:#X���0$6�r6.X.�S�q�o�e�����~6c_�oWSf�+j]AV���u�q8�1�A8z�ӟP��x�s�Rq��W$%�8��H��<���}ld��f�o$>�$4꽩U����\�&b�`�.zn�k������2��lS������.����Vʀ�k�Wx��>#%� 	�hĳh���`�Ymv\)4$��@�^���r�g��˗7��B~��=��Kxi;��U�����	|�[���(+�G�������Ќ(���R�"@��w�`i,��8���#��r�0�f4�G�w�qP�-�9�ű�Ǣ`k�v����SL �/	eJ���:
��ȕ���a��&�)VG�ܺ|'Mg(�N���/�3����bF�"4$��1�s~>�ޛz�@�t�1|jխh�,�.��&uhn3RHF�RPޜ4�8�3�X?U<�ҙ��EbI�L�ͨ�t�8) \�������_���A��'!^�=��ƮK��)�E��}vj�ѳ"5��~�eE���c�F��������w���d�"'7�2����7��5#�N'��6�I����fc#;��ߍ�y��ODB7�W���(j`1�y��]E����5��"��F5'���k!�_y���D�Y~�5=>��Z#���yz�_3�^�&�I��*�[��M�΍yk�>�:�5���3��� �!��"���Y��	�>,��=��c�"%��  �I��<�Lݚ+��� v��LCj�O��������K&�Q�FJ!\�{���ɺ�v��S�4~�:��'Ի��8z1��hY�m�Ե��<G�G݅ �qA	d_��h���bB!Ƞo�.�`c5�	���<������*��J�[?}{�V_[�"\.��9v�ɾ�6���IT�6ޫ).�dW~�B}��,97ty�W���iU���n��P�6�Ǥ�G֐��&BH�?���S���$x����mAi?�Y�~�n���xC�qg8�\���s~�_|�b�$�7�2��"��$l<P&�Zf��R{�RQc]2b{:΋�l4�ș�]��!�d�҉�q�u˚�� ޘV�IMQ�~V)�}�$@?I>t�0��������-B1q\w �ns���5b6ԉ
�}7o�mƖ�^S��Pd�.6H�<�P�ω�;��k<4�"ZM�+��\j�*�ȳ��+a{��SC*��0�?p@h�$I�a��wĥ��ha�L�`��:��ZF��uc�e�e�v!��wXM�$٫œZ�&A��Uu0���Y�럌�*����ia;��7O��nf���o�R��/?#
@*��~D�̐���ULfR����>4�F�z���(Ħ6\O�$���Ә4KY��|���2��}k<D��W�i ԍ�	� �W�e{�Ζ38�5DE�İx'ccy��Vͳv���<t4��(؉7�����w����+���sȻ6ܣRձ(�l�� �g42�M��"�����l�t��w}m�֦��w8��u�����}�A�X�aͲasNz�y �knl�n��V�O����
q�䮍�7ʟC?�N����ҁ��]��Y�4Wsp-2m��%OX���Q���,q3)\'�}\���A�&%�]^��jD��k�1�Ij���0����PګԒ�$UVH]R�/���-��
�Y��q��*E�㮹�m�_��u�s����$���!D+躁�S+��(d�!���:p�_3#�I��L�GÜɈQ�"�m.����Jp�z����j�&����KѤ�J�\R��
��L�+���GE���Z����r'e@W��T�r_㛷]D�ɴ���F���O��M~!z�]�^�񖆕o�j��\I����M�����<.�_Y;rU?���h���U��÷w:n� ����eVFSZ��~[�V�R߅`�;_�}A�D��~Y"#ft�b�����<(}˕�� ��Py�)hZ�kav�>ˌ�ys�}1ӧ��|�d��+U���.�Dȳs�Gxt��)�j��6�j�0��$T#v�Zb����}c�l2��������A�kR��S�I�,
(����	��8j`P�5ߒ���z+�f)��-X�*�hj��7@s�x�ca!c�rQ��$��� O�u�@��[����/|0��8����$�jJ�^����>�h	�f�*����ץ�.��Z�%�g���d�R���0/d����t[����N���O���u���ǄZ�Rc���h�m�9q��ׄdϿ4����WN�Ye����`=�"l�-��@�2��%_^�
U�uG��h�Q�YBw���¶cDgz�	��R�o��׊�@r�Hjq��A�uls�-ԧ(N9l���/�]"Ɋ9U�3�����X%�h��k�2=P-�����{X�t<	X�Q����A��h��f��m��v�(dq.Rx�{jV(hL��*۞�Fo���]Q����YР�[(y7�3gt�O�yN%��e�J�A��74�O�+�;�8gײ��_h��|�����7&<��J���x������j���ѯש��:���\7�U-h��n���Z����'�'Z�pA��y<s�]����8��#�o�.I������$jZ,M$�#�#�J�w�Љea������ Vc����ak������/?���QW�xe_�+}�[���%�`.6]�5�2_+�!x��Q^���i�u����f��O���ԅ��ѻ��k���u�p�W��\�B���A ��bn�C�.e���>a��b�4Ʉ��w�ck�.�o��A��=�s�
�4�{n�Zq�UCe�Ä�*]�kj��di�7ϯ� 6��ϸ��<e�ޢz�oC+��O�v�$z�=���,�>hͦ� �=��V82�Ev	0�^j4�ۆ)��L�j�[W#�	]튘���e�J���R�,�'�V�%~����%X���%ˉ�����_��\�'��Nn�_��w�E���Ƅ�]��_=bT�X��F�k/�6�gh�Js�xd-hb
�+�i�h��)3*I&���1�1�2��Ƃ��%no�f �sV�a��΀}������\�����z�d6Z����B'�x��*�e�E)�--H�� �k��j�A��W�������o0�+Ɇ��;|��2>^���X�O`���ze��T"�u����"���d��v53���@'��i�����U���NK�7ar^�-;!�~��KNK�ه����+��O/e�>�]ϼ������)6�ݹ��H�S����q(�sL:�	�P(}�|��KsA�_�	��Д��--sO�Ex<��������8�r?����18c���C!n��Z����Z뻨�o`^��m�����x�[^_���� !�N!i=��א�C�3hT��	��Yu���R5y�6����6g/
uˀVH�D�*,���A��6x��L�8/�MG��!3P�.~�5o�u}:L��TF��]���V�#6s������_�%\w�g<���7�����'t� �k4ޅ�$Ԣ +;����{ ��Z��FZ����;��&"і��[$��%^\��̲��S�V���G����G6
��ɩ�o�Im�(G��7m6>�G�|��k�#�AW#����cN䪭�n���1�εu�C��b�)_����2Г�/\�)ܚ�N��p��"hy�`��J�ů��A'jb�����Q�4Ђ�Q �Y=��6���T��a4��N��]�ɷ�Ԩ��9ٖ���j�d�G�:�=W�����W�7$�),�p��������9E��l�qq��P뵜�Nr*�����_��y��cz{l�ɗ�m]���!��m��w��K�����M��mlOG�D7���u�����~O�{����!5���Ad�������ʲ�	]��3z��(�R�����OlP�I���p�J�T>�m�?9@��L����6�IR_���Y�'�>��,�us�4k��<�i��]F���Y{����>N��I)�Qo<���e'�i���=���{�qs�īg�N� wtG[E�E�ݮ�A�>}^[�oHn~n6����{q��9ߠɕ@��[6��_����Z*&3{��:�&E�V}xjȀg1�}�[��n���!��u~�S�zq\��c{�=ϩ���?����K����VB�3�y5C 2��ͅ����m���d3�����'���׍B$8>� 2��3����Y�/^� �C�l�y06��x�&����>�L�G�H8�'^��T�_rw[���
b��Y���M��%�g�U��8;�u�$Y�8�Q�h����S���`*���<z�E�>I�sh�N�������sS;�]o�ݐ����4=�k�J���"u�q�[n��7�w��C��e9���~)�{���fD�D�4A��u�O(7��5��m�0n����rڞ�}o>��xY6Y�㸧z%�U1�8�_���iu�3Tg�`R�/��!eΔ<7�Ǝ�o^�+��YU��D+�4�;TY�:��J�QbN X�ύ��ZK�<��xY6���w*���UBqⷘB�uy�>�ua�D4���ZG�����v�uK��R�x��/QSv
]י3 U��<������G��j
C��/m��OTT^���R���%7���J/���7̹]!�^��G_��lS.���~�P�`���>f,hF-�"�K˩/����+��q �<����1@V��(s�<�Dm8~`-1�W�"�5qU���
���*�J����� �n@���i�ڦN7���$d��%�QfR \��C��A7�G�mhf���Naz�*fu���qY�n��,~�i9����%�\���|/�wc�h�v{��8�lI�|V3�B�at����η��J������<��#��0#��Hy�=��97�����M���M1�H�G��~]'}����;�}7���q�M�&/��Z�4�$�hC�t��� �rs0��u���p�v��&?}{�!k�R2u���֠����V$�G\�|�ee����5S��o�kRq�r�
,�=��ЅCt�r!St�U�.X�҇��c�Y�`�x%;�o��:�~>��@����ZO@�2���*e |�o���Wqt��	u����ߋ�B�9t�~7��
��>�
�PD0�h0FW$jq�᏿�f��l��R�')C�[�\�~H�ms>���D\For|�nͧl"�Q���,'�G/�\���άaB�d�������=�n�Vs�P�VF�p�:��S�ҵ\��y^U�f��sPrb�>-|.��JX�>T��[d��ł��n{}��xf��&������ugc,��Z��3���c<jWt6Y�qqĊE��s��N�S����=ѷP�pQe�IOm]�B߈yV��-[�E�@�
�ŸFE�6Bc������P��C�t`�/�6O�q�š��ł�`J�s�rg�
����z�QQ�!�stf��J�w���( �\Գ�5����Q2��^�����< ����N�b�������|e����[]��'�gl;�y<�*���,��(�b�ꥮ3�O�Y6#�O[lG4��4�\L,& l�=}E�xٟ'n8FC���O��ě�+
6� -��J��� }j4�c}�}J��� ++zo5�!��b��<�ؙ� �\剴����klP�/���b�� ���j}۶��dk$����%�`IL8(؃	f�kȘ5�}缨��m�e2�u7�����)#�F'�tzۆ��y�����;]���:�h�����9�Wb$vU��_s��U\i�^Z�\%^!V���h�b�dr{�Ȥa��_�3�v�4<Կ+�c�:60�1I�M������]��wN�Z�txw�����	̡�W3���tJh"�H��Ɏv�Q�F���Η�h�́�$��Xs��Kd�]M���@
,��=ڎX_;>��<[0�w�F����^H*�;5gs4��������w@x��Nn݇�E�v�c\�c�n@�`G�e^��[�Z���iL�5���^��_�`�0R��B5�-|��:A`���#<���+E[��t�1<;�Z-i������5j�8�����#ܸ��K��!�9~=Y�gf��4�.k/;'N��=�3_}����t��PUuB�)��H6��Vy���"}���E��=�j�>)��osRi4A�x��#�@%v�<J'F��9Q�����(�*G����v�س�Y+��Y��:���~8���pJ.���r�UR�M@2����=#�T��F���W����yM5T�-+Ug��d�J�h�W��X�ٝD���'Kv��-#���f�q����w�hyf�`����Q@�Y�����R��6�'��j�ᒌi�?Hf"|Z;���(� 5�*}����2�y�7�#��t�d��Y�K8������}- ���G<B�e�z69Y�`�O^�����{V���e���<=i��+��
���b�ϥw:ELJ�蓫�?vk�I��R����1� ��%����=���>Ki���d>�Ȳ�az���s�f%�#��#�o������HIr5�x且U�?D9���ѩݟ@i��_5Ĩ�2��ˮ3I߁�����b8����F���>=��$�hrt�n�L��0
�+U��U��0�f@���T�i;�;0�KŬs�Ȧ�*��~����3n5�>@4��I��'�K�����m����$+�x7Xn}��w[~���j�4	a��]�djy�t�D��+�����W?�����	�%��1J��t,c~m��V�y��ύ���?	"Q��%��e1��_²5���9D��)��<�@y���)����uB��<@�ǉO�cBu�s #�QZ�ŵ��R䤔���;mz�*|�j~��W���a|��,/3f��*�u͇���x��9^p��a�#ʞ�i�ԓ���H�彽�v�����Ίs0��L� /��9a]��mʇC���֙+A#�u��|�K���<������8�6ZiJN�N���Ɂ�&�gՉ�涣'wg�7���s��D~�o�)�&��T�c�ɕ���V�{�&�c��C��P=���Pf�4�
h����Q�цͰmj�T�y���9hVm�'}��>��&Ń]�ف��L�$�*S�'�6_2��w�F?�q�\�|�n��_m%{�|q�esSS=ޤ��5_�M쿓Qg�����&}[8���{fy�m� f,.D�l��>�P	�ҫ>����tv`����4|��020:!�s.��[
�(��U9�w�ڢ��#�LNsY�.AseG�����f� ��<h ��OY�U�7<�Է�5�;��� ,G�(Y�E��R��v��1ZA�m	w��G�R�j'3�Y�ၿ�Y�e�-@���_X�aI=᣼ۏ�֟)��"�0%4�7a���X��!zb�Bcu}$���e���މ~�#�����q�uO���>��Z̬�x �e)�)�ɜ���|� xdb�x��v�����ܳ��/n��̪�L�%�0L� c`�o�S"����z��ʙ���GH�uւ)j�Z�`Ne��>9�ϰN�a�V�\�]�\l��.`t�	xV�B@*ս*:�,&�$$�w���|a��w`>����h)�
��BO��O����M�	,U�\�=$��#�������F��M�F���q�I)�H=�oW�b��۞��9C,a�3�<K�NtGv�4> �q��W��ք6x�Ep�M������X�78�4	�V��ϲ����8b���B�U9�ⓇQ���9>"3��X܍�\�X|����GȜ&Hxڽ�SIE<#-���xj+K��4�QɿG�� 2�����[���ur� v��.��Et�����e�DQF���)��R�q��MKۃ��1��L�{�zyEZ[�n�ѴPk�*΁`�ɛZ)`�������o	�_Q�)��XO�<��ģxDf˵�d=D��HZ0Bmo\rO@jziH�~;�d|Ύy5�C��o!8��  ��,�
ފ���X۲�!K���Kt,��ŬD`%�=�Q���=�X(���EŚ ^��%����Oy)�7����l�5g�1S��~�5[��n��ڌ;�J_�O�A��V�� ���<�而��������b�ި�ĵj��y�ÀI[D���z6�lih�v���W;w�vi��1��3!�ɺ���eH�W�����mW|�+m�. ��!ۼ��߸y M��^Q�w�/�O2����z����Ś�G�)��L�aO�!b@u�v�����S�t|H�9qB���ߪ����c�}�g �0'4��*|�ZB�ʦ�
>��J�.���a�]E�9q� ��f�O�&��E��M#4�,�����M+�)��$z��w�+|&�LhGJ>7зja�n�q���l*oܐܺ��t�s�8W�U�C��
����3\�F��p�I�$u��,���fr����t��7��%͉�nq��Nt�]7H����H�P�L������.�1(�.��'��XL�婩{��ڬ�T���_	X{gD�ɸD�5��y���+ˉׇ!���Jr~�yw8�N,���j���w��`��J��sY�[��Pt�3#�_H�^��J����BQ��3���_��=GŊ��RǼ���`7�|��pJ�� ����9d��7���U#���^�6�͓cO��rႶ���?K*rX�4�lԹ�,ģv�Ý��go����WYS.o�X�L�����\�fn�����:�<} �Mw��������!��U�+sܶ'�Y�"�Շ��-�k�US�,v�Fav���#W�Q���v��5��\��'r����&�	���M�����V_�i�5��Oӟ�OI������I��-�X*Nr\~\�7�5�UB��xd�ՙ��l�8�u
�W��rB_k�Ds<-#�����H+o:��L�"�n���ڍ�o��`�Jz6�Vgm���6b�^m��ھ��v)�^��߉�?5�`�/���Z�6�qL� ��+#;��B���H���5�Y���K��ѹ]���dq�-���4� d�i9z���()薸!l=��׵�E�@P��-fQj� ����]f[�j;��)A�Op�������!;'/b�KG��4O;J��R{Nf]�<H��:ዅ{�X���{ι��H�1���"8�K�U�l��0�k)����t��ҭ�ב7��z@���l�?Y��Z�IEM��<��CC�n��1��)�E��L���s���k�[{�
�n���������1Z�rZh����O�u5#��A�J
A�@N�Wuv�C?����=mz%kF��{��iZ9VW͠�G��9w��rg��<8 �ں2��K����w#H}�R��J����'w� �ɬ���@��ւ���E2��ϭq@/�J��x%��&q����.mg��[�A��O�A��T#o�v��B�9Ƃ,�R������!{�q�c�T@(0\-���^d�/� �94ҽR�����c�7��X���eظ�/�	�#Q�3,�&��2w�F�{ȴcyW�����C�7h���+yM���r]ȸ���n�p�q��@Y��u6&���t�hݚ������ [�R�ֵ �6��_p�רk��JG�C��a@�W���pr#�p�T�j��Tyb:�R��."(h��]"�[(��h��C��p��w!�f�ר%�����y��
���q�����/��F @��k�����x������k�i�r��Y�y��c<���d�Hj������������6��"���`�F�x�S�J�����A3��X��BꈃCB�ic<�,�U"m ���eԨ;T����8T�n��!�]:0c������~|Z�]�F|�$�.� ).��>z{'#%(P���>\���7|���T��Z2L��59�ϩ��a]W��6x1���hS���u�!njR�#�;h��|H��/�
�}���� >��7[��2E�E�����V,;q����veB�Æ2�6l�(|�J�Y��!�g���J)d�!n�Y�YZ��6�h��I#�ͭT�1B���{�vc�qO:��>���O�� 0�c�2�y��x4��A(�Uo"Y�uT&��Kז�JP����!������ ��C��ޒ�S� ��#�;�Ea�]�I����aɤ�|�/m���I8�Y�/�6��f�D�(ЮqMM!��Z�ޯ0�\;U�0�ZPJC���uU�D�>Q�;5��^�����0>	�@�v����%9�}S��/ނ.�|�EY}�����ӗ`���O�0(!G+|�1���ߖn{O֍��߶g|/��W��|��H�_eSs��vep���k���кZ��?�l���v�+ݏ"�(��{l��shub�g�t=�� ����e*�uR;�@7i�p|&�?\�a�t����cƗ081k�cw����C.K8m�V�X/w����k�B��Z�r�#)���?����/�j���E�W��I���l@32����_��qr�ʝ��xkgH�n罵�� �s� 7+x�}���E�lħ�gLeDII��r��P`�ɞ��w�W�~�7 ���µ���<����Ϲw�t\�����k:C,s�;)��2�ʙ���k�`�����
�eJpˇ�ؐ�Ӯ,���QoY��G�D<�MFEM'Sr�t�&�c�r���������V�A�a���h�]� �{����&j%U�Uj�p�������Q��:e1ǚ�������n��?X�/"k��5҃�����/�i}�񞼊�P���^E��H8�3��W0�k*.VK�/���V��%F~�+�ëU�<v���|�j��)���Sݛ:�r��ܤ��p��P̏o=�ў��'��6�ы]O��2�9=t��
;���zNK�ay���\S]�A �L�s�<�d����-�<P�VFY�«����	����(�]BY�m�𦢪k	dA�!��/�u�n�?�v/�k/r�xTT�庈��B�9�JU92ٹ�fΕ�(w2J�7�}��+���(6R=%��jDJ�SW��0�����'�"�]�q��U�X�0�i�q�9<���F�Մ�#^��1u����:�j5n�d�Ƃ��� ֟����R�ع��o����SN��[���η�Qar� ������~�QĖO�����҃������R4@�[���L��5̘nj9:�D�'Kͥ�3�[�Iq�^�B:�O}��ġ�am)($�6��^��: �6Ϯ!��,��fr:�����W*=�W�R�5��F�Ė�F#5�YW����5��m �W,��n"��xv��O7�����%��m�z�:
�m�d�%����|;�@��{izvf�ի�EA�r��,;��eU�;�Q��,��\�hFɮaWu����X��Pz!�)��M�̧�P�'#��ó�������~�{��׸��yH�щ�=4���RP�Q�8e�vXmHk9<�-2������pq�'q��-d�e��떎p�k	����R���~���t�u�����O��H��o�)�ZN��{'bH�u�g�8�}Wa�zÙy*3yk��Y
x�q�W��"��q��6�R�l꯷�Ԅn������o�Wܪx�����1g���L��m�"56�a)]pHǍYd���1�:��8�ToF���h��p]ϝ��h�M�X�?6<�u�p���	�-�/�ls*�9)8�������P��l�HaHא�Ѽ4/��K�ڢ�VL���(��]%e�{v��p>emy#@���)�����ʚX����0����X�!Lf�����\�v�sT�}�p�2ʥ�l��FĊQb�W�)rµ��h�����3^�%���b�з��K��Ng�/�QD�\ !��Ɯ؉�Ϡ��O���_����$H�9���xTps��^�~ES6Ѝ����oj���B6������]���6Nh����L0��A�x��d����ަ���+.�sO��c�V�N5�k�	����P&K	z�m�b�	p��Ϻ�؃u�u���f(A�j��������gh��zM��q��)����s)���k�����<®-Z���L�����8�omTL��ݟk��9�+���K��k� �)��x(��}�{��[�=<
])��Uk���/"q���zF���zȑ�H����ڴ� I�/�/�)K�1zĢs�>}#��!�� g��ifV��a��9�pjȊ�E	NS�A]�=ny�����CC
嗵����;w��o�0���R�8�t����^=�0,�J�L�
*�@hf�ȏ|@P���O�2t�U
B�����)H��|D`fO��h-⒓p���ڟ(�}�b�#T�Y��iN����d���Q�$�P*E�:��n=�4<<-,��P#1Q/Mn�o����R(џ����9>�<�J�	eq���a�>w'��А���;Q�Wu|ș�J�/���"�U�2ӽH�Y��on��W�eQFǃ��d9�}ѱR�\�^�l.Ȟ�O�;�Z�`�Z�(<��� ?����|�#�OƇ��b�k
�]��K^{v_�r)j�l���I�d�$�	��߾=V{��Q�q����uPx=�0L�ɏ8���W#�7P,�0L���fۤSE��i�@����!�	2%���#|���F��S7�K��XE��g��0��LZ]H���5�n�7��蕽]��5!�#�6G���7Ϝ�1�IE�y��@`�+�O�}ӅD�v:���;�ܲW��� ;��i�4�H��M��-x�i5HǕd��t��:G�db�/���ߵj��	�^X�;D�[ҝ�G�t�9�1�1�M�)�zAq.46�5q��]<'���5uٱq��v�8�V��
l>_�%(Y��e�yւ��!�KZ�\)�g3�$4�I���[��$>K,o䙴�e�e���4��2f�l��
�Kٚ��;���n��n��ȵE��&�&�P�.N:�����rc`��ɐsֈ��)�Y����0�q��U��]*a�
^��:t��_�&x��Q��E\��_�N����zoa���.���ƹ�O;|���#�u�w%שW��J��!w۷�/�,|�
{����(�w:����]pk��_s��^�i����������P�7ӏV3�g��Srj��3�R�Tl�8��'�ӛ�5�C�A���u���F��	�ɠ8�;�vz�\;Es�i�I�g�?�dxi������?�#���m��Ӡ�!��C�6<Xf]���
�Y�=D�����G���t�A�[��J�"epY-�l����yg�KE��S�z�dy�/1nn,
�VW�S�N�I�SA]e��}b�����. �gT)��������ē�:L��`�l����ž`h��`�v.����2n����1��Ћ2�\�Φ��4�14�
��&\��U��O����_�8a���m�)�!�fi�h�+�U�w��4��÷u%^eo�E��B������M��gREN������])25oT�5�G&-e�s�_�iJǾ\6�eݎ�	{Pܨ�͹<>��6Ej
��#f���au���W2�j[�3��ydۀ�H�R�2�;��4�)4+�0���QS��/���8�7� ͈�VB�$O,J�P�����Ȗ�Dc�}�F�IQ�l�X�O���s�WV��k��yL��_�7�P���ny�d�����J�Xe_��er�����kaJ�Y9�/��G��NvM.T0�	�"R��uT�Vdp=�6���wl~�ZuҘ�&LBc�&��t��<+
$<����I5��&��|�/�̥a���R\��B
�qr1Ȭ֏Y��Q� �ꗮ��_�f��KH����`�Vy#J��j��hI02Cڗք�>}n����+�@tw0��L�l3b�@�-l�=�#?�J�Q��ܛ�|������Ҭ}x�a��W���m�"�f/��}[I@o�����%�>�쥹�gt����� ����žW��O;aJ���p.A�0���3,��0@��@G����T�/ev,��AȺ�T���7�$`=ɉ�_-	��샚�K@VsD<b �[j�o����	��M���МS ��w��O�L5�v����K��0|>M�����NT�_�K���	mWe>�=Xxf.��XXw@l�����1�� [�cKgg�̻`Jg1�w_��%1�����HouՁ����B-'.��T�A(&ďol��3v�ճ��A|��2���;�}� b��%Me|M�E�j#�6��cLmԗ��Z��T�1���T,y��P_��d��4HW(���V���r�Nь7��������c����-tYh�eÙ�۹�+�i�SXS��m)h��ЯAg�f���ףF6�Fv+rw|�V�l�am����9/��zW*pG�o��`Xp;�rK�-�5���!R|V����C�'VS��,��a���Z�=\�eV��H�=�׳�4�9���IQ�݅�hZ��b]!��� z�;��?ƚ���L��˛�ΗJ��'"�?�D_S#��A0�%�� ��|�PwM �sÀ�v����;��/�WT�9��ͥ��#�k�LX��k�� �C��lo��:w67��4z��s�N��Y��<�������=��s��Kx4�bN�T�c��9`�:m�K��h�3���z�@P�J��Luy��u)���LEƥ�|��fV��5Wp����y�y�������!^b���G���R�����:�o�c��e~v�^����B' D��]Q����N�XT"s�Yp&ۆ�X��,�1<�Y|�qF�Tɉ�u�-�H��b7Wя�F��LV�z�@�|��e��`]p�x���b���S`�W�6��cBd�x���s)]޺�W������*����FXJv��/����A7�pN�:j�AA�"�c�q� bP ��v4��1��b�b�ʯ�9�f����<��:�y�6Ɨ[��':�S (�0��~!n�ب�p�x�l�����nP{sp����H0���@oi�c�V֡0r��x����Ç�5�:�.�X�C�:.�uK�n��=Y���͕zg���8����U���e�����_i[�|Z���=����E}��pD�0Ԉ}m���e���fJҦ�o_���:�E���<!�a��r�]�K] .�gp[Em��D �P҉�ưNɈ�w#E��0@@�(`�t4�c�j, ����=�v��YW�H�`>o�
�L�#�!2HV���J�8c����>�;�������c���dZKZK�q�=v�ۛF�<����̭]�ϖ��L2.t�
8��Px�!�c��R�PN��nL�H3s���&2�Qn&Mnp��Y��{tU{D�¼Z v��$x�s>L� ��JIN��XZ?!CQ��ǩ��7���k�M|�� ���C��4Z�ɏ%�=ժ�ݯ=����~���+l�ř�4�Rlh������07`̈́�M��9��t�[h�� �����y����
5�n�{�L�_�(�n���rT���_�i���Sf�K���ΪX��u��HW��4g��D�%�ܨJ#֌|�گ�v�fk��|����I�BǼ�[�2�\0		ϵ=l!�B��w}E��+Q��b��ݶ�i�ME�<�KP,s,���m�Z�) w_�%���kt[���IƎ1ђ(H ��Q���/w�VT!5j o_hJuw)X0�"�ڹ���>%@��B/m�a|k}�;t��� ��=�|8��ZɈ�:�1�%�����H���\��'ӑ�©�j�Us��E�P�e��v��"*���O0P�iN�����R��](��j��zD�$���d�)��X*�ﾁ q�z��䴸JEH�idn�i;mt<���d��>��Σ�� �� �)��iI`�;�?���0W��fv��3s�_d��e��dE諺y��Ή���ǈй#����n�n��#<���-OfGc���N`�Jx�F~7��WV���^���v�~}�b�q�.���M�q��鐓�� ��ȹ_�wr�\x�4UQDFyGa��O���<�~*E<:9�5eP�Q��ӑ#��j��N�T}��c�(�=����"m�|�7���{PFrJ
�{�%�Zs�	�&%�fN�������nb��b��2�u�`01]5�ÿ/�Ӣ�zVT����]p���+��|*+�EH���}*�&�)y��i�V�[Bfvl�6�mB��K��V��TEYc�U�oo�o�:�[���a�[O�	]I�ȟ��Y�~<xQnp�K� �z�w[gq�n�X�_^֫�V\�\E�^�G�8�M�x+��a�GF�'����SP�C`�����]C�����z�������T U��K_�f���wM@�I���0c�igF+�t��<�7A\ܣ�!+ܘ�����4_��2
�R��q�6(k:6"]�\��@�Xd��Yջ�D��Ճ����n\��hN�����K����۲����&>lݛ��<�R�2hu�3Ԝѿ�����vN����kD����fF�N����U�l���C��	�������N�� ��f�Ӥʂ��`���� ��>Z�'�M[�@�X`�KT6�����}gV_@�Ĝ�f�?]��m���n��HHXpQ�@�Ӊ�5[�5����l/�wI�&A���y���~M����#'Fz���~����6c.l���:����U����x�Ĥ�H�x@��}�t�:�(���3))��	У�=H�⤝^���~�M���N�Y��s���Q&���*d�B��5�\+Z�P��X������s�ӏ�c�A1!����1�1�OA������)�GME��ǯ���߆��Wt}`����� ��-g��Ұp�)+F�%3��.S�q/Ł�J�Ƿ��-�P� ]�����rw�۳d��B;)p����_�����p��+�$X|����Z�F�e��F%,ڗ[��_��Ryd�]񍡩 ���'��կE���Y^ۋ�^�l�|0���>;���a�����m+4��錭�g���RQ�H!�����E��rb�t�>��b��̖3���gI� ~�-!;"��Y��?��\�`v/�`̄=di���h�{e�5D,����Q��Z���u ����k����o(��]x��`����j��V�!�Z���ꧺfl�m�J�ZSGV?�"P�]����q�C�[�Ө5P�N_w��c	6@$�g$:��6�p�pP�/�;ka���Dr�/p1//�(׊�J��|�h��#���3D���J�RP����0'39�T�檫ޒa]*��<M�W�݀$$���l���6ȄH��$��<T��GX�:�̡���[�o�];"�&v�{��e�y�չn�K4��#=<D(������w6o[�8�A�A4�6�(e`~(	�l\|��w��S/�2��	�!v������	���(�@.���˙��$��>�Ⱦ�2w	�C��wW4�9n���@��Ʈ��}E��nǵ{y�]B����
w�2���!�E��5%l�ܳO(���ۺ=�$ �V�'�Cx��R��C�O��+|��^Y�ш�������n=$�}fOf����=K�d�$�y�l�d�<��B�"�9+�j)'T�cL���"oiC�,�s���{=�ܫ��A��r���.ʅ3��qX��]r�f��7�X�4�@Ԛn���9?C?8�Ϸt01T�B���39�X����J�>q,�ol8K�����������㖾sJ��,��XK�N�w��A�;v�=��y�����)ǖU���Ǎ�A�~Fh;*U��h5�o�tm�''zs�[>�msL�qN�-�5,�]a�. ���Di���0�����	�(d|!�O�7<�+y]yːe�o�v�*��
��L��Ə]{�V1	��$~\Œ@gdz1�ӽ`�79t	�1?6�����$�_І��ϟ���R��#i�����r>�Y�O1���1��x	a�{c��c͕o����'_ʿfO��wGy�M�>R�)C�`VG�����N�O$��;��ҹE�  P¬H�Q]J�G�|&��rZ~����6����	���v������y|�@Կ����?U�Q���?��� � 7���b8 F�+�9!}�,8�M3e��|��va�lcx��'9�ze-Es��-�R�@;��Pލ�V�=����ϸ������ W@�K����Z�qW���T~��'X 0bwHv�F��{���Ì�����U� fR��2=�b7=wIw=�r�3XbN 9�x{�Fۓ.������檵��(�nS쉱p�}��&�7.U����C�o�/�W�{�ZK�	_������`�?V)2u�&�y2�^C^�`��|z�\�xǹǔ�ޡq�gQ2�L&��WN�U>���mP&7����/C�YJ ���X��|��.[�a�=�����a��|�>L�9f�?'b^�^hL�7S�י�ޟ�w���i�z���:	Ku�]N��G���-�
dKG�vB`�<#����A�F�V&�ݳ�}C\˿Y�D������ͩ;�I���8�5_�(�L��~��s����ݏ��{�k �]�� L����|��`��-��|�ng%d�T8���}��F!���%�8�!)�b;�� �Sf�f<	����,`OQ«�/��3{f�EER��X�����kdg����$h�g"6Oh�Ck=]�7�q:��ħ���}���B�}��{�-�+�(a�b�g���;��� �2�C=ŖI���P�g����-�m?oÕպ� |S�i)�6������|2�ۥ�ԫ7
���� g�7�����?�����*ρ�����7t_�v[f2<��t�!��t ��r��uc8�fYR\
�ef��Բ��V#�Z��o�>��fٍ\>��7({�����'@��J�Aw1єѢD,��MQ���ܮ5�.�!:Φ\8��|!q��"f��o��0�L�A����	i/�����oҡN@u��`��m̈́k��X�`I�T�`��,����`��3��<x�9�_� � ��N���%��x�L$bivS�����5*d��&�M睺Z��{�f.x2�!D9����B�����Rz�L� �O���o�������E�"<��ǈ(Y��?e��y݂��o
"�`�7G��:/tN���l�^dWu���F߫K�(āSEؕ�ب��Gb}{G��wkT��ga�x+����i+�<�t�l7�/x��ת�Xr;�ҋ1�����|؍�"v�bv�<��~�!e�? [�z�؄�g֊�x�Ա����6�S���R�	1+��C��"]�-5�ւ�:l0��Yk~��1ͩC|
Ԫۖe����a�����2֡R��.P56/�S�Ņ3�e05���d���ݴ�L_�o���xgt�JI+(��D�j�4�3g��rA�=��zs5g�|�o]�HV�$�5P�H�E��yK��#��� J)�x�,�g�m�5d57@[t�e��r{�.��4��
�x�uFI���x�׀^/��&Vݳ�V+�x�7 �m�f�'ޥ�&��*��V�_��i�G�zI��ɣ��!������-d����������bVl_TN�
}?�?�D���/4�=lJְE ��S�٘b*J�=��P�)j����g�%鸫#���v���G����M�A�~�W����#���W)�Q�Y���*��5�SI�x1e1���1�:ޮl�`ƀ�@���+�����&��>����N������JkP�f�L&#����2J���A�'�n�I�A�;5��C�if)���$SӼ*m-��:���# d&������g�V.�����6�%������س�9�#��.���ȷeq^l���-F��ޱ�͞�&AO>�k�s%���3;� Š���pR��}���FA�.���T��_%n	�z��r��C�
RW�=Ǳ�E���j�����������2;ku`�%��]���{s�.��(������4��D���B�X枭0>�4A������6;	��<�\7��eDT�'�X��
޹�Zĭ��ӳ���8�������z"��"����̈��Q47]�5V�V
��v�Dc�\R�'�-ơ�2M$/>���q�����e  }C$_{uhdd���MY��xQ�i
o,��8��p��=^+�1E�����Dz��z�b�t�d��	�\:' ���E��5�1�yEtZEOUx�Y
���[�%���hxr��S�g9U��� A����W�]V-�Z��l��S�a��
��<R6�;Q�5��3,l�}����Z��Mg���?�[Bfo8��l��:Q7�iηM��Ż�6��0\�<�>ww֕�H�Dq�x�ϟ�SB�V�ɰ��-�U�X�|���å����)�΄�Kܪ{��c�BwI�]�t!TJ�k���f��ԎA�@�E]h(8�n��oA"�@;��|% HT��kE�=����R�B4���o��E?�x��_����8�Oo ��`a�Gച��)mk��/�\��:gk���W���ր/!?�A8�M���
�9YP�����Y�V]�~�D��n%I��Zy݅�u$�<���g��?�ι�`	yP����م�N�e22$x��t����g�܉����i�xr��a���V,��=�59�\��;?G�8��!o@��UA˗K��'�.���=y'�
R&�'�B���\>�m��ڬ����:w��W�j���s�O��+�}�����U������"��G{��Vlշ��"樯����nSJ��S��~\T5H@#�L����f�V8���IbiG��ع �Qe����Pz�оX0�0	$I����yY�5IC���N���ofx�V����0���1����b ���X)�g]q%AW��5+G^=L����\ꈴ&���9~�&����Hm��G8\6�3Z�]3כּ _M̔8`i�M���RY9�9Q"+�����>�ܒ5���%�#kS�f�`5]Z�9���/8���g%Җ%�z�8U��^x;��E��l��z�'י꽤ؕ�b��&%�$��rI�5ܹ1 ��|�� ���j4B.�Gc����L��e+�@�S�YA�W�0rQ��K�G*�ƭ��a�z�E�̏��g7�8--%&M6���f"�W�^A��/��\��$�.��(���=9�_�-������N�܇F���!uq<fd�W�H�䥝9����Ƥ�8�&�r��G}.
��!��{��W���b@�ti��n��+��8�T��[@���cDZ��2�>��l��֗�d��he8��@5h�Wʡ�e�������<gn��֩��Yw�	j�g����Ǧ�1�lh���Kj�K�h8%����:4�+{^M��T�hFs�W�ت�&V�3`�o��)A�A�i��HI����r!c)���9�l�.B��F�L�UM ^7bnA���2�RwH�6Y��\��֜D��onȒ�b	��ΙJ6��ԵAU��,b��Jˀ���s�}g�vqO��&--`�'Pqt�HW'W�CV�?;vͅ	dn5���7Z�h��?SB�V�>#y���b2T䆜�#l�I�0�#�$�.��0P0-ޑ]
�6�����vDk�G���'��%}�3���|5��#�KK���k('���]�P��n���Ω>�����BS�R�E�Q�X6��'�1��q�CQ�^�E(Q�B�3������ʊ�O�滀MZ��u�IF?��W��6��&}��q�)�wR\ ���u��ldLw뜃��wk�=���d��c�!��,�N�Q��!t�9��!�+v����;L�\J��C�@B1H��ϔ/$�j�g��S����f��s*�Rm�������̍����V�ͱ`�G�}u'e�.F2M*t�U��srɢ)^={7*,�u�sVnd�M��ᔐ��y��'���+Old&�KoR�PC�/L��,ۗ,�yg)�m]��f(,����\�P�N~F����B���zDLՠ���������v�ৰ�����+[�Z�V�7��N�߲/&~�����'x!�aO�w4��W�E�sMaa�8����X��& �R�|5�t"ؐ1RS�/0iL���CX:���#;������� 1v�p�E�JqMyN0��]	��"i��ޜ5nw��`����E�ꆀ�Z�/R��(ۻ���I�b-�<�������cH�ZjO ��?���J���c�ݛ+D�����P��d���8ˍ<A��0�l@�{�� /�q�^�૮�
CXql��	U�"����>�P\�����6-�
FF<L�j]T�8�B��4_s=�*�/��fd�c�u7��(�(�G6�o }#z� (nw�b!%Y�@H$��B��y���8S�;�1�<���|�����*_�fgH�鎤������㰜��� ��
�*�_��^�$U�k�j����l����H8�n{���8b;3%�F�}M+_M��r�K�Ev&������cѢ*h�Jv��	L�wOI�6��V��H�WYZ"�4�)`�a���T�;���@\�c3�&���t�CӋA7�ݰ�S-� xj ~au�& ́����N2�1\:mϒsDS�.;X��/�������ɱh���Ŀ�;�o��/��cK���@C����*�n�_��r�B15�Uj��S�_ܙ�-��:��T��)���@�х-�c�6N��V����޻�zt����D�0�Ŋr>Gn����`�Yv�Z^ĉe�T�I>$$R�E�zTI�iqZn �$��z�����G�"�-]�\�4��_����O(�-{�O����}�J������퐣�����@3:6��|N_�UL�]�.�$�s�.D���qN��a}�(�q}��ɣT٣�S�]�:�̰VXcX��:��w<�a'�w��T������� �3�����7#'K�k) ��Ғ�;bSk���`��'����"��)��X*�.�6ʢ(���H��:]�YXHۜp�o�����2�ު���>\�t��aq�����h�A�X��	�;�3���_p9��t2Gm2)NiE�~�/8"C5¤��l�C0C�<Pl��H<[�"pZ������Ms=Q��G��"NK.�M?o&R�9㬠�w��/�V#dcU�T���7~@^�I)�r{p@ƨFU��� m��&�1"��pBg�<~2�2C���!U���tl�v�[�q4N*f���^l/;Kp��_�3��V޹S	��S���91[: ��|J��E����,S���)^�6Qn2嘨�@Q � �I��9�K�9�np���`q 3����P�f�4����4�<Cw��[H����\��븯&+,�A׾� cvf=zMҫ�(��@�='c�60�E=87�#o7������f���ۧ4'�؆�M�X����v|��� �D_��zU/�����-TѲC�I�6�p������O3e�/��K��%Y�{+�~��Q�l�m؈�qφ���t�pg��xV�]k�S��&ed���֖(S����듐�s)O!��|�l�nBVj ��D^Q����3��6`v�<��Dh�7!/��j����"����@4��t][	�"0<��3���/����	c5���ԬN��(��o�5 VL��8�}[4�|G]l�;��K'���ٟ��+$TEw��������I�~���㊾u�G��1��5�T�0�h����2�1�"zO�a������KB'�����]ِ�>uUT��K?I��N��`�֝�s�~u�F�v�;��	�ְc��dt��@,~c9����飼�g6L?Ķ���1ڲ����w��l���
������P���h�6�L�B�4+�Y5{r.�}s�� 3+B9���Q��L�߫�����V�Ip�O�
������#�l�N|�8����4�!�M���>^N��!���P��"&<��<)���%մ�y��D�g�A� �sHĴF�n�̱Lm70����ń�ҽ�Ν[TL�Rp*��5Z�ɏ��s"3/�=l��␎2?sۭ�묀�TjL �H�ǿ�x�:a�4Vް�$�TL�[�U��G���>���ԋYo�-hx�td�G�;�Z%%��`&��S��酑;��o#y�D,�Km֊�+�j�]�]P3��7�S����Q������h��wY��ju��=�U��A�9�c��΁��p?�Py�H:���a9(x�hRY���g$�;!]��F�_,���N0�� 	@[��Ʈ	�+���vId0L�����4{C�i�lr�v��F/�+	"�l �mBOg0�f�R.��xy��_���F��zt4'"�|6$���U����۵��>\��&��0 �i�X`���y��
�$ڍ��؛Ⱥ���n{%����������'I�����7��������;��Z�}��Un*��v}\>��\���S�L��(�R���xpb+�g?���{�����{s�sv�z|�0Vp�̐�	�#o�J���.!|w!��a�Z��s�:r�Ѝ��;	�,xnHJvQ8����WN�%���*�V��|�W�� 넛�	ԁo>�����h�q�l8�FԪe���"xi��a��pΙ�]����JNc��n禯a6R����_�#��{�s*�hÕ����e�B���?y��ʾ��U�;چ&�^��W�j���U�����ޮM���`�}w��3�-􄳐W[�2�J����ΐ����.����Gd��=����Q���L?���*5ʻ�������p���� d�g3�N�TGUy[�.�q�ܒ�ƅ�3�{��'=3��n�����TK>�R�xf�L{�I��Ǧw*�^�G�L�UF���EƔ���}@�F� $�y���8.!J����hU���U��q�)S {�p�h��+�jsI7`J^r1�I�q'�6��Ǉ A6�"T��G�"%���[�|�8K�����E�j��ͿL��O��e^ci�M`V��(x}��.�[�KR��A��*0}&ʥk����r��" �J��&1>�ݥz��Qn���)��WH�%{8]z�	Zw�������C�ьW���K|�ϰ�(�a>b�N.J�D�,���[��*5��kik'p� ��g�ٯX�޷�7��i���x��9�.� )�nC�Q����C���0�*} �]e��X]G�DK9�&�2��Í��x�xM�%-�#��vL'b��ð���0y�#���=���;�R�VX���s�+Dd����$�Z6:ُ|ʝ�����.�%5m_h[p2��}�d�oV�w����e�{�sO�i�G�x@YMw��9|��o����9 ގ�o�����P������"�P�?*=��!X� �2�%�,J;�E�?��ŋ�=��P��!|����6�?�\�E��Q7`���RQ���A���wd��[(w�%��y���,[�_���M6e�K�s�f�X��oh@u5����D�G��ذR �Z�D�4�傭�G�$�#hhs���*^D:�x���f����/�'A��VK����֝Y{bXɨ��ޘ��!�R��/��&��ǹ���^�'�{;3����MyÿH�Ʌ�V���P��.⏾��P�����,�lm��L���82�& ���6_όa �R("o�d!�[ �]�!s���G�+�*��2^3�i��c&���XϖE=��=���1���!I���I�����ci��z3w4o�6�������
��w`�b���n��˸#��':uX{��ō����8G�c)�����W��dt8	��{��{��%��8����B]���Y!"T�D;����te����,c���3��Ȥ���J� +��W/�xH�s�Hu�E�=K8w`�	+�MZElT�;5����C���Ȫ!�������c���F '(������y����s-p�W &�g5������0����	��������2%��tn���(4uR�%�E�Է�Ph_���`����|�_,�"Ө��^�)|m�3$$M������c�:�b�H@�2�< >�"B�����/�D���4���i����h�tw7�S2��BoW^�T��m��8]�k�{�\����)��,�G��.k�AD�.�r�M����#���rK���d��JrY;I�Q=�L�+<S�T��4{VR�����q]���QO���Є���c��M���?�0�:�kI�OU8��2�Շ�Noen� �{�������"/����;`�̔õE�]?���,o�V�+J0^��ָ)B\�~�����Փ�80.�O᭳��%*7�[���8q�����2��9j��L��R���k�%��q�+Es��8(�)�E�3OA�Qci*��^��Z�e[��GV��f&,��g/;_D����1��bR���W��<�`�˖U�J�����?�7�sy�*l� *���sx�/���M>):�|N��O����o�m��MZ�a<޽�?ޖǓ�����ts�c�u
�u�r����������C.b�h��,�Fr[iW&���~�0��c��)�e����Z�'O\�~BsAM>4,�^U�|oG�e;�;�;��.	����͆�!�H�l�H"�O�]č2;����QŨL?��@?;-�m��{��}�aM܇�:3���DS�C݊�M� �k`࡝�����)�AS�v��S�S���g�I�B�JG%�d�|X��ZZ�1�{/䀔"�K<i���֨�����5x	2�_6�t�I��-�J�D�?��!ܰ&�ShL���;2�'�o�I=Oa���v�!�l�.�ӎ��Uav>a�2zW���͒ 5����,{��&�;qAk��g���-Lc����6�I���+9�a[���������k�>@WŴ�l����q5��$�^O���6�`�� ��6�k�s�̆�������kk�_�z{S�g�^�JvM
�ӹh �{��1v�-9}ʧ�b�ȃ�Z3�������,?���ak�R�!�C�����6_�_��l�Æu�M5�Qΰ��۷�v��q�����ȓ�����c1l�L�*��U?TV�:kxe�5xP��EPHw�!y�Jr#�M���ߛi�(���	ps/�~Mѥ�&$vS�k9�c�ʚש��b�},:��;�/mΝU�����ME��l1��Z�K;+��髐�����ȠjO��"�	���w�n7�����L����-�#V^����\����C�'e�bZ�a��������H�/��5,��)��#qy_q��+(H��M�7��-�����<��U�zQeVdOƴ�!݄���0e���{�#�~��pB�i1r���F������?����o�9�;�&e��9���I!�fj�<��QPh�����b��H1K��HR���<�����g��}�=O��x�,�f�/�( �!��eI��	��쭮E3I��I�L��n���PU���_�ˮw�����smp����o�ֻ�kt�`� �������ފc�{����"C���^̇���Xua�"��I>LX*F�-J#�1��dC���"�y���s�
��l��Z�o���z��2�I<wj�Np��X��e��u|�_qR��O��P�v9�^[���~��� (���̆)�1�3�v��#��v}$�/�|���o۪����<�O�f)�g)`�|;Ө+��0Dŀ�z?W+I:�Q��fK���ACNs�#Κ����/�Q<�J�n��Mv�L/Q�vb�\���i1��k�����8m$�
�y�=�D]:�yP��3�3��<���{	�6�xS���B����t����*��8>�(1�[�=1��.�읛��BL�CM��nY��<s?��_P�@�A	�	Q6xJ O2�J��Q@��k�b�@����o��Ws%��U�F��ev5k���T�m7V�F)�=��\��N?m�ե��!S^��v�V�0K;�ԥ�!8U���9h �uz��ٳ�w�X�x���E�
��<��g��J�{�F̟�st��#��Պ#hE��c��5��m��uG�C�d�Sڴ#�QM1��歒18r�ԕ�J�+�	� �]��Z� ��i�h�V�s�L��G���H��%Ź�2�#�1}�����ڼȹH�=��� ,j���Q�w�����d�uK"��*��;�a�)��E�����.{7X?_�Q��0�A� ���I�/Q ��Tm��-0O�W������?��;��*�T�2�58���u�SY�!{S��>�2���{]�g�?~����P=�m[����m�G�\' U5��������)ԧ�]�!B�4�����3�$�(������0M��`��)�t2,�<���ȷ%O}\�rH�v$Zs̊'j��&�9���-�>dn�I5������+�|���I��zօdF!�0��{X^$���٨�3m�by	g��w�f�O�٥
q'�x�bJ!]�%��Q�NwlF�s�4�}A1���7���r��;ɫ���6��?�)��Ux���D~t����8O �����U��(�)��سҌ��qhRV8��k�K
�^o�C:��&ţ���J�`VK���y�k�y}*ݨ���@~ [LM��W�|��p���q������U>����$�G�;_1��u����>w�T^�`�����jE�TPt���C�tJ#�yӈx�ڰV�֖s��]�c�������g������%���ƿSy;L��VHS+�(88㟀�}֒�4��o̖����Z)9��R��۞%q~Ɖ�g,�0݉���/M�7��fhQ!��l��?@߶��9�t(e����dR���K8/*�@���1e�2��K�c7x��zN��w�Ϣ�X�A�G3�n���;�y�؋��g'�8�\}�B�ET&8�V�/�w��=�^�ƴI{�r?^�x�V��QJ��k������-�-��ciM{m{�.�֗�=[V;�0����}#�nS~��1'v��Bl��!$b�l�PCJ ��u�>�B�{u�q�mS���JD�*h��-��$�	a`�G��M�hJ�(e���Q��g�����Pd�Ҷ���A��D\o��~i+���Qr��:�{�H��``	=�~��{����d��X��ݕBqt(C����6�r�	K��)y)�t-0�	6 �D�ُ��߶��D�@6���j��ψd��WF��ѣ�#�`__��w�5�̩Iz�)���8�0-�.���0%�m�k���J���46�}��Ao��jN�TwPr����C�6/��s��S^̎݋�Ƌ1v]2��4��K����7s��-���
�K��w�>䔡��"t��=&�1�rH���C}���,�ϻ�z����3={�ᖛ�3u�a��*^U��}���R��>ȿ0T|�(��L��@A�B��:����L���Gq'��-@j�g;DCC��o�\p^��A�P��*�|S[=J�4vQ���9R�u9͢�E�°PZ*\�" ��z\DsoA�+W'�x��G_�S�����8�fw�z��;͢* �щ7�M�Bc�Y�K��8^Xљu�ލ�����uA�3�}��bj��2���ɼiG���\�Y�1?�-��~�3P�җ��G�	\Ҽ�ݟ@/u��n��GΎm��-(��g�^�_ ���0B.9V}4 l��"��#b6���2ULgַ�I2�Ws	{~ǅ�H@7��۲��/3����,�(�O�����Lх0����%�E��(��.]f�E/S�5L�C���2�
g �W�"��.�O�ݓ��s���g�~�,�_���8�wBq\g"�p�e�&a��9�,���4WQ���8xS<9�ݱ}r��l"j͗S����8�:_�	o���G��� ���kM��u�=Y�- aK�g�,�Q��wu��|�`Y�z��N1Pw�8� G2�W'�o�.�4w[~M�A7��eĄ���`�Q�� Oy}��q��c��C`�g`YU#�vG�Tw��S��,�u�p��mo1N�zy㋯a�iEK��2���A���%��]uj>�ȜTZ���[²��6�,*�#�8��>�ߎ�t*I��"�|��4��  ��'�A+r"�
�Q�R�=LO�IҰz����w��a�S�q-�+n$�q�9�������_�[�"�X
U�[�����?߸��Vѷ��'�%��q�ʟ��w�Em�61�״�0J�2D��p|�'���~aQ�]XTK i()��(�s&���%f���t]������~���aăf&̛\��(E�� �Y�G���B�L����	{�b���.��=Q�]A�C#��IT��|]A�w��Í���9d61�QO2�cΖ�
��U���q��S����vsU��1����S^�|�><���MVefט'��y�L�:����g��E$�~o�݇���A�+X�k0��6Ot5���F��sʾ�G�e���O���̢W��Swq/ژ�~�bh@�x �.��"�E����W`y�}�+�`�D���A����߈L��e}�3�+�!�_���ek���^45�eAf�0MI�Y�Bd6�"�ፘ��������˹��&]r�	IG}�6��O��%��"�oXo�� ��'4��ʗ��-8�5s��)�j�wX
0�'X���B�BgS�V����N���͒�� ��Ͻ��7I�Ik��%�A�7�w�����B�0h��������S=��8TM&�֛[T���E�z7G<r��]��bҩjS�NZC�	y����S4H����$��  73j�jZ��(��<��).��C�me�Cb�h�a����ƴ��j�Q�h������B� ��ڝ9�5��[x�;t��mޜM���D�����fQ_�	��G|ƈq�MZ';cp��w��B��E�~�ˤ/*��p� �a����؜���Z�uH�'�Ї^D �z�h���.)���;���
u���#��X�ﻯ���^ʯ��9ߗ��[��"��'"�)bH#2s�h.�6��ޛ�H�+�]��R��9s��TdO�H(�)�G_f�����m�#�E<OSCa��f��E��m]��i��4�7R�tpe�'Y~�wl�ӇX�y�O�ϭV,�*����P���78ֻ�P~OU�*..��9I�Y����9�p�Wl�����˿����C�zN3S�G'����u,�'�2�0��9.9���I��@R�N=Y�q���]	�qZ�BQe[-��I~�ŷ6��e��eFD�cv�6`G]�0sҷ���c��0�͑�����3!���9(��I�m�jVPDY ���a�	� ÆOkJN��X�3�䛼����e�i�cu���ƞ��uF�s+%��]-�������F��w��,"��%%�b�wd��[��Sc�#m�AL)�c͐ª��>A�īA�\�n�Qԩf�����Y�ͩp�� ���l�h��M�B�a���A8J��)�T�6��^�JUO1�S�A7X�{�G�4S)73 -E�C�2)�Ay�,��w���d�2��a����u1�X��4�-fu���l�S��aW����фQ�Q���"�@����%�7�k}S�
cD��}P��*Q�Dn�w�i��$"{U�K�Hy�gS��O2�A�����F 9�Wu���M��e-��,��5�c[_H�6�͆ۇ;^v��԰:%Gc���~���8�k>x3��1<aW�����I��P�R��J(�0�s׹+�h��ѕ&��9�����&,}�j���k2��dC>��4K桹�S`��t��e�O��hr*��x��S\W��<Ld�t/��[� �gxuY�M�,M��s�Y��P�
h��A\��8^��+�*�r��w����	{���������H@��Zk|Z�&���q<�p�ͫ ��G���pP��&S��zHI�r�Ww'�=
T�I��*�?�0�(K$����pd7�i�e�v�#�Ɔ�|��{b@�54����5H���<��䭺�No����nx��/&
Z'��B7變i�
�2,'�.�9�F-���&|(:7�-Z|�,t.�Z���Yh^�\��CM����W�p;QVPN9H� e��LK�}o�W�G���,݄M�u��I��"p��b�_1A���g�������eOm
<�ɍsE��SX����O��i��~�5B��^f�=�ݾ��H��{]����U{J~ʖ^�틻��o2�
W'>��	�5�-T��r����Lك��ͅM�s����b�����]�m����d�Ʒ���V�:ln���?�ՐW�"b��8n/����DK7ՂR�L�c
d�`�d��L�}�EpT T����I��N�?LoZĜ.	��E���<^/gC_a�%�FD�"�	�PK�th��,��8z��׌�����v_�ք D������:�%*�V�#��_�btc��T�y��&.o�����idg�5	b�At֟���nٟ~�����{�m�:6	�(���,�0�l�X�p�3�r��^|I��� ��X�k-����m֍����c���'}�x���V����ԔEl9e����K���swu�������uѴ�@9��@�D�ļ_�!�D� *��C�$��Wj���*^�ei!�Io{�4�غQ�n�7����5��,���|ᐱY����ô!�M'c�憆����3���W�o�(I�]��$�,���������<�[��Ҏ���LUV��C���A>u��+=A��1!S\�ɀ^wt��_y$�=����-�s'O$��Bܻ�{r�_���S�o�<����Ե�/&N�#���{��2EyqD��9=#����Y}F(�"��,�k����3�����u�5�7�u�����uF�`���)��l�T,�"em:��{vƙu����ߡ$�N�f��a\�U��֜y�89�yg�mYzYq�L�2���E�:�"k�P��q<���ENЪ�G�� �M>�V��e�d"vX�;��N�6D�����J�4�<[��x�����9�q���H�۪����nN�CT�4�8�C�_�c����Zd�b��[���\af��f��K� w�p�G�-���}4e�ڦF������Q1`��v�,�2E򦛫��2�枠*Vr�������r�s�!=�𠺓�͙w����(�p�V�!P��>����9@��Xͯ�	���%��Ή����o�ڃ�fp�~�q6VA��%#�[�[/����`3����R�t!�|h��F���,,��`�����n�5��WۏyW
J<�� �V�f^�YT4I�_o�;b927!��&C#�����f�͓�T� 5�Kϓ$��(������
q��
��y��/�h1�;x���ԠJ	.S&�=9��Y��H"�^u0U~�h����*ۑؖ�a-`����u>]��9�r&��Px��V�<Ҭ�\�hx6�:/�=���He��dF������F=�+%p����ikq��Ck�r��i�Ĵ㙣)^��#�d`Ѭ]W��9���|������0��o�.0����#%�<p�k��T�����|��@�c���EϚ���RQ�@��
�b�>�QP�!��y�뜂)�rWG��ma*l��e򣙡���r�7 �5�R��%"]s��J��R��&Ҷ[�ֶ��T&W�Ú��y����|���Z;h��C��<���e6��������F�������P���<_��A�� �P���8�t�Za�$�"Y�˒���a��v�0����m�	��k���Q$�j10��S�c҅�P�>�!���Q�����Ak���?٠،�lXT��>M���:Y���5����ĕ�Ukx���ӷ�����d��U��u2l���\UJ�s�Ǯ�#!1)m�5LM�\�^���s5h��y�r�>m����,!����%�;?�f�Q6N�]����[2�O?�'t���$G�䠂.�)Y𧮱!+$e_j�)!8�[,�����P�xd�(����}��Ұm�>,�y��O��|U�s�:�Ee��!���I�T�� �,���)��8���u%^��Jz��[x��A�*������M�ߐ=��d�ӊ��;q���+���tT+�Bp���h�c;1F:xM��-_�3�,\��V��Q(}7�3ܳ��t���W�\ ̳��Z��������1��@��a�:��SU���k'$��ߓ�I%���?]���r1�甃�/��I�I�i�Y������	���7%�B�qp�R��#����AJ��A�%W�MN���QL�M�O�$�u�dzW��{�: cS_�K��4x_n��L?'
�!����s]D�.j��5�&�Y>%s�W�:����~�'�F3 �}99�ţL,��X�c1��[�E8�=ԙ�q�����[�s��;��N��1�C=p:T��,鬞����� H˝|�,����;2��3w��7����$�.�cF��-�`��>$���2����_Z��h��1Яwa3$c�A��^���f�����S�i!o�2��n�/�&ௗ�S�����H�N���
����k��&Hz�qK?��f�����~x}!�"�p�wBJ{� �TOՊ��< Cy�~XW�vCU�������������G��ۺ,1���XԈ~��,P�JC;{ii�'�Ԟ6���@?�K��/�r ��5�v�p�Rf�ܟ.��)�@���ēX�fH���� |��g����&~��Uc_�:���0�Q��B^��1@7�~_���"�.y�!����B�Iw/}r�[ f!�>����0�6��ly�#�=��D��忖<�{p���},d$�5�gsx�f�+C�a�v:ziDM�����Xʏ��g7�O健���UgI/PJ�B�&�P*�a�]��~�7�8S�x�{^�q]#b�l�?f
�+(D�U����#�-�f��9�Ysg끑�ݠ��` ����i�u�������:5� ���W��t ���3Ba���*�w���>[�(��z��WO��(PPU�/��ݜ�'R�-�[����/�BL�.�#�v����`7{c��o�5>�_��E����(B���Xg�z:�-�V˒��3��.�,<[%,�#YG�Z�b<�	��%�ΞM M�mL@�5�1V��$5n8�IĐ}W�RA"�l�8;K(@&	���R)�R��?#����/�Q8B{+@"��]v�L[���D]��T��9��R� <���6ݖl������9|����l�-�J�ɛ���7%�%�y����{G�Y���Byx߾Юj��+��C���UHJr.t��.'R����<1UP'��"�Y��U͍�˱o�8�V��+����#X���<h�����~��?�����"8�����TÜ�ݦ� spl{Ce0f�}��@�˨p|�����O� �(^�eS��V��E���\�x/��|y��Wtt��w|q)\�Ϗ\�Gu����$::�������q�ץ�1����x,���J�
e�Sm}���08�=P߃���i�b���^"�l5gzG�&�ܖGW�@٬�wy��:�o3]qcV.��L��k�n=`�����w��:�(�P�/�Pg�G'T�2���Z�[�7����������4$�>%X��#�+�9����]lz~@m��ծ	:��g�w�0$�d��o�/SR"��()I��K�o�[PI��1�h�wfx��ԃ	e�?Q�AD��խc[�1c;JΔ��m��Ajf_��c�U�P#����N+�vYl��6F�~ꊍ��*�>�Uy�5�(.*J_C���>%7�s�Z9��,���{��YZ潃�2�:��#}���&�+�6ؠ��"n�A��9_V��Bh[����Rl�*���m���*\Yq�4X�RN �B�H�AI��n���{ �具�+�|.$����	���%[�uoa������n�C�`xi�!��I�a��D0y��8�S�eCHl#�w�T���F�t�&DC$A���u��m��)��Ϲ]�X���H}ګm�X��%ɂ���8QB�s��0Rir��%U@{Cu$�kb�{��8\�����r���ci����O�'��3O6���}�l|
�@Z��=���Y�d�J�	x\���fɢ����v�o,��Ш;��!�̢]�X�W�~��f��Kjכ1.A�8�y�/�ǧ�,PpIҘ��h������i RKv�`[y,t�О�QU����ro�� ��tB�A�<=�V��P�r%����_k�ְ�	��͖ƕ���#�&�iT��m3�++m�N�ʨVӇ��7��fnO�-/`��)<wd���j�+��g�=��pn)��-��݌Gn��Ş������-*FX;A+(�`Hƶ�.+�H�G��]v�l����v]��{zv��I�!�J���$�/��ym��?2��P�n+l}x��:aY-�C�w��"�e
4�K�i��D���e-[���v(��L���ǆpMy_�R�kDT�Mڊ�}�"{��X_��e�%6J�7X��z�?[�։���ک%f$���5b{n��W���
 �ǥ���1KZ��Ð׵~Oh��m�8�T��]WH2Aľ�v���[و���dY�2c��]�sL�K:��1Q����7�_�����@����Rr�I�R` V�u̟9�jaKː��(�r<�I�b��F�5m�͌���7�	�S7��,*zx��_IO��&^	� y#�.��P�����/}��Y�O�q��m�[�f�G->J������X�g��f�<#ddh�1����ʌDm�����+��_�3�'�V�	)�1
�Ua�YC���h������y�P'�������]b�mt섛L���?Ʋ�.���������}���X�Ƥn��{ہ(�	��ǽ��@|����}K������r]B�h�� @|�	z��(���u�e]1��g7~���zg���O��w�Q�^���X���ڐ;����;W�Q/�*�DJiϡ�޷����ˉ�Rmj`*z���:�2����s�vn^eY�ڣ�Z��s�9_�p`<��I��.�e傭3v�3}���`�+���|�q�hQ�A0���bZ��P�EH���u�g�]w��U0�;j�}Sϋ�����pb����:sϒ~C�j��J�D�m�04��B�3�2�p��,����@)T`!��h�fG���[#�C'�~�c��%���!O[�'������" G�(�X:P�jN�<�
��z�ë��`;�M&���S�v���:��'�qL�FF���M�%�9S;�D.6=f�\o|��!�`d
�n��k���f���Z&Pq�t��j1����r�B,At�|b|j��R���q��oW�փ$���%�過�xU�e4����Áo2К��ӟ�v�CS�5�p#�g��hZ���|�{���[�@�����
?b���v�����';��R�������U�d��l��c��j��;����el�)]��<�C�nf��}�?oFr�ϣ�p�����
R�Fo��+m�P�2I���m �ǟ*"Va'M3c&��<�IS��`�d[����n����QgY-CR������[d�6Qr���m����A�K�
�o�������	-y�w�a9�[Sh� ��!*�7k�����ki���k��E�[(�y�N��cq�e���W�����p�HH�{5���F�@<��O媄+�?���=���H��9G
�
ie_�x��]���{#�@rh��X�S�la�(Ԓ�U�:<Hy��j+�&��O��+�u �KZ�yc�`��j�AbH����&R���)~����B�Hv$�va�)s�)���ֱ��r�=�ʿ��ֵ~��A��F�ūO����T��q4T�Zˎ[$G�or�@�>�X���?�}�G��F%9�T�;�Fl�nh����@kO�]�t�o|�X�}��o�?X����#]�n��Hm�!/5�{��C�\�>0�j,�Ǹl5��:�(�����8�%�RMfU����W=�_ZI9V�w���/�������̜����g&�9����,�����v���ބ�c�H[�a��KF傒�Ϧz��"\"1�7I�Ш��Q����^T섐c�d*C�SN&��!z���4�8�d����?�lL��`�e�����j0�=�-��&�	�F��Z�nJ�Kv%Zy���3�"�ޯ*�i�@M�h��e���y�t�ъ��A��~G--�,X��5/^�*���r\t�#�S��?�x���R�72����3Cb�D)��7�	

L0���7��'�hv��g��u:H07�l�͙@�{��#�B�Q>.�c�qD���;@��ۦ�D���2^1�\ц�c�I7.H�����#)� e�iڟż.�ǜs���?������/��-e�'}j"��N��:6�{�����Txj��^���Q-WJ(�E�j��[����"%��+N�����K? �?�S�2��?X$�4t-�����W6�P���% O
+�3U�d8�R�q��}�m�9Ӿtcwal�6 �������)��{���8�7�a���ld���W���rNͷ8�������Db$�s8iU��#p���LgU�  �t�*Q[�_?#'a:�,c�g^>�]Rg29��^��l���L�������B��(�-����h�}$���ց���"��G+aal�'�E�=�=�Yh~6F]��ҬfC��u�.��Ņ�N�LT�C���K�/ñ�����桊q��zB��9��0nbK�7N2��c�]2��N�ɀFH�EI!�%�k˷S���_بSʹ	��u�R��f��u�B�D�@��������j�i��9u��Z�T?�����d�� .B�1�]�oT�ٷ3ɄH!h����[����hv�ؕtv&��UW@&v�����u�0$ȟdj6��J�#��$��}����:�#ŉ�Z�=�����W311���k���
�Į2���Wr�pt]^��siV��va�+�(�~�g���;�=?�^q�-��f4���4l[��L]��o����x��]%�3���zh?�P�:/�!J�T�f��g�s2=6�t� ,�s ]�M�u��c9��J�oWW��U��r&�hg��? ;�Ǝ��G� �XX���N�n�$�� B��7�%�Z�eE�[9���l9�M���������s����{3��V���g��$\�"n��؝������-�,���l�o_��6 B.�6/�^�@�a��i�d=;�NZX�Ŏ$�ݟ@��e��Y�--�ײJRe���0t��*�l��5~�ze��K��u�����-��5�u�-(8a��a:���$n\���A��dv.�o���!CV"�;ci�"��5��Y��݈� #�h���-���o��nY6���h6�|�]�P�v"xJA�qm�ؠ4(�R��R�"�w���+]��j	��������x�J��n]1XDd�$s:���KrW:MV<'�p&�ܷ�����F-�Q����o��ҏpn� 4�=�W������)	�Wx3��x��U��4~h�5Ew�ofQ���?�a����2� �.!�C1�^��L�e�X���rE�4�o8}��:w �C��#�ּ<��Vu<d�d�d��aZ_�5G!�� w�|]�U��6^E��"v��u�tf?U|7��	E��N��kng!{�07'�'�����JGd\�]@��#���x��[�ԒU�[Bd@���[>��R���Z�ޅ������0�k%���s��O�����G��*/{�Y�k �`C�矗������sEy=���)�����a:�hX�� 	�4�i���q�7%��CSf>�?��6�%u;�	o3B��2��������<>:�ρ=r�.dYk�-�����Xޔ['��:0C�Z��	��r۲�T�|�ڏ ����ޖ�ucY����+f�K��}NV��&���&CO�1��� ]y�?^�� ����7��g2�Un���?�>�k�)�5:h��Vv�*s���k�p%-�J�mM,��Q��e�Y���Ό�G�ZeS�f�ě���S�v����/�G��j�Z���x��a�9��p����9�vSp�4�M��2��6M��Wgf���0X��
ʢ�1$��ph��Y�&���]�����#J�͂B$P;]�qI<Ϥ�f���p���s	֋G��b�9q�~~��%>7N�G��v�n���"L>gmQ���c�/9Ԟ��r�7�%w�QaT0 �9h��(���߶��=��h���ϾU�pCF!���6a	�/�b�B�`���������^zpe�S?!'���!+��(�G�u;ٹ���AP�SI�����ʄ�{�=�hs� `�c4�m���������]�8� x��I�߶^�������g\�.��\^�l����u*~-x�Ȓ~�e��h��9Yw���=`t[����8
�~I(Et,n���"X:>�ipe��%>˃%2hR��
At�A��T�y�/�yw3��6�_C��IjS��ʰ�KfG��!��^,�[��N�
&(}%�jL=v����w����ŶZ�_;fؤ	��+vG��të}X���OF��8{y:5��k<Y�������`I�$*}�X��۲��B�^�6�R�p����~��G"E�g��P���A�tu��]L�6����?o#�?��n�?��~^��x�����:��I�����{��xi����6@����(W����"Nn[��]  ��µCK�EKM��D�־ݯ���e��*2�'e�y�;��%I?�| _ѷ�O�XB	�=����'k����Tq�<=��.м����Ly���;�7g6�p�[��+��l��,�������S�{.�B��hz	@G�C��D�q�⽾��G���r�ɧ�����������>1ђ7���Q�nMXk����L|^��m���V����{���d�B	�͢LZ��DĪ�ʥ�DV#�Lg��c�/��^&�d�{�G:ݾ�sm�G�����qU�Ja������_����i~�v"l��aN��O`^�m��#2��a�f�X�}	�Ps�d��H��0��R�z�g���5�J�U����<2""Zy��R=nAAP��e�C	�&�1���
f�{w$�h�	GMTF����K�|��=��A��<�%"�⽰�I�l�qK�<��.�Ƽ�7}:8� T��`,<���@���οpW���xf*i���@�h�%���l���V
0��>��91�*�����L��A��7�;LK�`����VY�G:�ɶ���8�1�p��%l �eϗjy�&�OR�O�}CO���������{H�J�ug��CUU9Gro����`<�!E�,*�K��0A�0�m5��"#U��P���h�M{���e��0���XR�
?� 3�ۣ��0���,I����q�:���{d^��'	��3W����^t=�L�]�׾e��(����eU�#�����P�|��x���x�j��cdU=.�H%��snb��x��3�B�g�/8�k��s�G��=�8�	����_j��Y�#�q��r�?�5ZWI6�����/�w��v��"�H*F�X"��@4MwcCPi&��y�`(^%ch��y��7��&���V�BHQ܁0�D]K� �G�Z�I���T���i`tO�ͥ�k
ٔ!�/����D�Ƅ�Ej7��@�t4����G���彶�خC4
�[�
�� �ʛ�}lW��}B����8�2m�% �H��IkΫ^?��u�.6/܀#D��'���h臺�j �..ҺOu�;��h��n��V��Y`��,}&k"%z���MF�{$��<�=#�m���v�3vA.=�iK��<kJ���x�Z�&�5z0�ŉnѓ��=�Q=�e�&EA�@)y �D"��D����1�.=����(�5i�}[J1��iߎ��v7�[T�%�)��4-/dD�F�#s)���t������b�F)Y�e��C�W]�<(o�}U�, �z�MK x��k�ϻ"A�k:���a܄:,�k�V(9��:c|i蝿L\��/=|%�T�o~]� |����h,�ͼ~Uu���f�82(��ڹò�!Y��f��ЭX
�.� �jc��C�|y�@�jD�ZD��ǲ�y4�����감�D��C�����K�ĩ��Wr���]@���^ ��p��@y4��Qϝ}��@|���e3���5r�5�tPN������M���\	��A��.�������-SV���gw�Q�!�Nփc\��*!�q�q�wM��s���;���͆!�$�V��I>���S�_0k�[�r��\˩92�_��� u������;ͣ��`�d��P"�֘A+��Y�����<x|Y�A�VU��oA��+yČ�e-:��Y�G3��C�0V���k�rC�a�4.i���� �����G�p2�B�V�4�g��R�H�;�S����wJ��1�u�O��S����.M����@�b�P��.d���Y�	�9�ZZ�n�I����&I���TF�I��=]�GZ�B
��S4�ɑ�p�]�F'�=��ef�q[�
������s�ｗ���	W݈bǶJ�U���6�QF�t?�ft��B�f�H]1	��>ćBI����g�Z��q`B>$ �a�D�DX�T��e�ˀb�R���#��D17:Ѡ��Uz�CT���g���Ca}{����S7�)��} g����r���_��Lh+YC&�8v1���αN�;}�Ό�EG��]���S��35���g��XA5܂=n�\�ˬ�.`E�.�HָĞ�k�f-b0���)\`���w��}[�����N�Ag�H�%kS�. �da��ёD�+���M{�<�"߲�o�V��J�$E��l��2��Y�l���g����G�1{y,��1�@�����Z-n_m��pz�>�k�� r�cS�c4�������m�E�Y3�/+�KYs@r�A�G/��Xy������#����c���X���9�?�������AcP��y�Ѣ�tc����钁|�H���r/o�ː���$"8x�˄��oHH/^���������``�{n��Qm���dc�7Ŕ<�.����cV�o�����V��6�p%��QR�C�[���T�aD������>X����k,���6+=�x����I29H����JxW��mM�WFj�ߵ��S|�m�Ŏ��yh!E]�vb�N8�|�B���U-�"U�����hǸ���Q�FL������6t���=�tkHo�1��~�bb%3Ο��Ŝ�TM��?(�%�W*}�;O\�2q[&	�œĉZ'��OD�*��
�=j�x��H?F ��L�$h���9k�$�Go?]u,���DGm�4�$7����մ�YյF�U�;�H��/T�1|��i�y�r������	Ν8��[M77�G������;��3��;΁3`/=�Ɔ�e,t���![[D��C˙���Lwq���0���F��Կ�k1��B�'�d�T�[§�0�������D� �V2R���H�|���%�����Ho��鲗�P��D�E�	�(.�H���v��p+z&7�"Y�o<�nr��ᭀJT JH?�������������a���S���V�n)�&���xN v[)S�T���SmXr4��@�\�Z)Y��K�Sc�4�L�)t��{A�4�?��e!½5]��o�<��I��S��t*m>š����?c�cU��/ ʇ���-l`�h������V�3o3�qڲ����L&o<�~�3Kb��*	9�ΫrL��G����K~a\H��~�m�0�Ü��^<IV
�0�o%W�PB�5�p��&y͙L��!@����/���ͭ��ԙ�s.ϙ�3�v�I�wC`pv�ڔ)�D��/��C�g�g���E��x�!��3C�Š4SB�S��i5!��B����m8���f����}e��_â�<�������fn�=���h�q˧��L`�f�\�>5"���I�y�u���`��SJl��=���Fy>x��-���sԨ/��n.�Zɻn�jYH�@�,�ߤ-����Uci�#D�Sh�7�f��s뵷�^ E"%�g�����{�7nu�`�O��4{��Xv������{*R#�gc���8D�g�AOxͪ˿sh~M�~�q<�ԑ�=V�-�F��F��4%p��Z���Z��g� l�U�u��xLY�}mb����>��+��j�7Xy�H'�CF�ܦ!ԏ���������B��m6�Ur�㳃�aݔsˇ^�M�-�+�ƻ�y��k |U��׃�gê� 
�d1��b@��ɷ��I��M'��;��lGy�_0�F��T�t�ս�~�n��}����v��4�tH�O)��� �fe��G~w�ٲ�I���*�®4�h٪bv�)�2&�&Wj�%�&�����Y��1��C�ג�=A��(8
��@��m�9��\�ſ�2"\��\D�Ɨ7�C�L�[S�i�مA�a7	l�t�"=r?Go*s���h@
�_ 5n�nS+�d48�H���amʀ�T	�V,�Y�ן��_��/Q��8�݅lb���ΝO˖�1�/]}|JT�����~4S� %�s�J
��q����P�?}�q�]���*<���Z���a�k�u��*��T�n�I��\)�+�8�"V�h�.�j����'�������i�FT8�9��сSQr�I�&���>����_�&���ҿ�Ӡ�]��0�u(��7�_�W�4?�ό�9>N���0+�p]��"�!�~[�[�W��P���n�j2�G D�� �:��n��
R~*�8J#�MU�w�m�������/�ugK�q���g��]97�1t>j's��D�r��肒_H��ɼ��J\@�W���`��䣓t�;���]I�t�{捸x�� :��h9�_y&h�+^^B�⊴��ʝ�{�ta�u�ӣ=�Ŀ���5�r4�Q~���q. �aC,3ͥ�5�\��41�D9��=I����}`?�v��?!b��&Nt�0QfP������7&�S�m��Ӹ�)oF����KG�#��U�e�+�H�S���P���ב8��T���O5	)֛��(_�1�7ZL{Q�0����ؑ&p5���0)�����$�����}�L����-C�H���3h=��ǈ���|#�=�VjE�������NN@����ij���9	���i��4���ZX��+��s�������e>8�i��|�3ٗ�5�؂]�����j��\!6r�����O�X/ �q�*;��Y�������!�%̲�=����G#I�LW��b��ھ(ǴaRb�`4A
�Q����)/|������@���N�^hm�2{�ˁ��h�R�W&k� �h�xd�5R1P��R)
$:�ypѺ���D�v=?FWF��|�Ɔ�M���P)wa�Y؞�P �-���Rm�q	��gk�W%�0�2Y^(BTB��J��-�1V��(p�,�=�ϴ`�5����hAX��d`kQ�L36�� o%��9d���.�e.v��ͰQ�P�����=����'��8<�� �BB�.�3Z����Q��7>k���W 7;ُ��,�Yv�[�`oAУ-9�4���.�	E?s��sR�\��|��޾L^���T�Bv�60B^:��I	��%x&�$��$�Ŝp��LW=����Xʑ���sm�^��U�i������X��,T���KU����~�B�/M�c�b-��K g�ю#M<J�$�����N�Q>ox��s���&��Y��8�-m2j�V��v��{���;�a���ֱ�@{K.��M2�?hJ�]���~��e���aN�o�ܜƔA I�Rq���$�J��(D�@�~7��m�hg�:B_�aL�Ѷ8<��M�X�H��h��S���
>xL#�Jˋ�*^D{� ��R���H��
=-���O˫��������~�D��2:�_���J�&q@a����W�F.�?�ŀ�[17<(����?�JK�Ǻ=��ݫrw����DrVp�kmX��(�(����6��ˠ��z��#�`���΂���{1o�-@<	�LΛ�?t'֗l<�t�t�M'*�hF;6��!}��nG\-P�V@p&T�`8߰�֜¸un��txUw��4������q�.�e�0�<p|?��P�e7�Fl.P���ѥ��Y���e��GƵ�u��~:F��I�6L�~ܞ�p�-x����h��}�yV�jV2�(�&b0,м����@ſ����I�j11�R�#����zG��=b�Y.������*�����"8�!�<��<^�@1�*�Ee)�65룶"#�cs��']1�{Q����+P+��z,�g�}�{�c�E�a�L��%hXI�}u��h�"�J0��-�����-D�U4�`C��;.M��{�6��Ɯbs�0����I"���D�S�nCaj����K+w\N:�%����Ƥ����Mױ��1�� i}`ӌ����G�ؓ��(7s�=�H��F�j\���_W�dH�
bE狍ÐH�d:�W�N;�Z���vg��ݎ��|�[�� ����c�M�T(��_:ߺE�13�{?T^4�B�Ƃ.i�Z>rt��9q�Ũ��I�N9?�,�dr�|�������h�V��Շ���T�R�+f��ɸ.i���	�h������}��m7��,��+��:���}>��,�[o��Й�8�G�4���D�g{�qY$a�^��\P�ŒTU��E+��A�v|��׃��^��2C�˧G �"8��Z��H���漋C�';jW[|e�afJ�U�lt��?�=�(�*����j�k!J)�xl=*��'@����s��5r/���C�#u�^�nUY�H�������kv�k�m�E�
���� .�M~����lד~osNO��f��Zѳ�����ɪRr¼��'@z�Bp
[�+���� �&0+��Y���7jٍ�c?x�(�q|�8!J�C�p�Ȍ�
�Ӂ�>��^@���9)��o� 3�\�k6A�m%�$�b��A��{�c ?�p���"h�D=��N�*��][�Ț/�Bc?�kam��Y��L�Rg�}��I<a~�Ċ�J�_�,��h	���� ��cE����Q@�nJ�~s�2%��Y�aJIM��i0�/-�HS�����AB�T�Ivg@#��'�-�SYwڊ��z�w�!o�I�KW��1�k΄��'Z�~=���|�T����vֹ�����V�9�z�DơS_6��"Z��P�ҏ��0m�m�I�ۅ5�a%�i�]�G��[���~��>��O�2ݑ�m��Ş��a*�_�!���1l9���`h�S��u�7
'�p��Ƕ�hP�v')[�`����+Tx�7��'<�D�f�I؁����p�~���|Sin���{�]�M�A�u�߈�C�p�td(��&:������j0���w;�0xVj����E��0{�c����HF��8�7�˄֭�-��v'F�� ��t�����Bi��ע|:�$��}�JU�y��4��Y�Km�:F,�[�P�K���1�eT���/�@�/�� �f�s�
����12�ڰ����$Q��cD1��E,2
�3��]�?��KU�?�Bd4��RwJ�%�Yj��j@#����F�c���ݚ�i؛/�����t�W�@ܿl
��Uf;z�\���5}Հ�g�ǒ�-�1J�0��[@ ��Q�}���*�]�E�
ɖ/���������t�F���BU���%5
npd8@-ǌ���y�$���b��6q�t��m������i� �;Vx��Lr�o�^^���DC�;����"�]	#o��#ZZ���c�X�9�������`r�����E�(���񭂘��hGߧ��Y��4�ah埕y^r+�$%����Y��I甋S�Q}����{���|�VZ}�
ѐۈ�6"�kK��7c�-�9��{��|KZB��b��x��i8.��$#f���H�ۀ#C�����i�"'ԫ�p�$;�ּ���16އ�u$,r�B�
,'�8�Y;|30j�fG�Y��F�8�j�iDb�6i�3�^E1z��O���<����������e4�T���샺=5R�Ǚ��2?�I�����׽��iIJ�5�͞ʒ����G�wQ�ɴ���8B?^[�5D��f�J&�3�Ry�X.Z���V�w�D���|l'��	�󊾦��V!��ha˄t�p���V�-*1�}���=����a�m��&Z�)'~�V�|�R[��խL܈��]¯��6X�O�8Ie�p�!���Ö!-�D%o�œ�#R !	�#�x`�DZV`�&o����FF펚G_��߈B�q�&�C�০%k�$���ծ���J�Ǖ�q�D.�r������?H�s{�Vh���0��<�!�EP
�S��T�pu��-�ߤ ��cƋyϾ��hp2ñ�j�j��@щ��k����7����1શP��nN�C	��U�7���B��0(q|S��7�g��hx�$�;Y�r�$�e��avݘ���0�Ƹ1(�!V��@�^;Ҹ,rp��3 �yD�>f�SK���D+�f����GG�?W��!�nF���˱��l�K�O]	��tGGO�s�ڬ�����%�^��W�2��Q��;c��`9BЖ
�9�m�i�R5탦��~$���N(��Z9���bB������|Q?+'�D�E&�+�6�[`�){7���,����γ�8�lL>EK�`O~�a�w~{��E|	�� ��	<�-7*�&��j>9|�{����'/-�$u��^�ƨZ�Ǒ��ޟ��K��ݵí�Lq�H,+C�Db��4�6�Y����U�M��!t!�~��3V�Fݷ�	�3�F�A��F4�~��j����	I���`���Y�s�ן�]���P�h�GY/X�"n��I����d^�+��V�An�K��:�'\���]�h�Y�d��qq�p�S��EuA��C��9y�ܪ�Zun����0�=|_h��OϗQH(���ցĹ�=�R���\v`Z30̋#O�{'N�+N7��.4uѬh)�H�z��
�<�v�ж>�����6�����C��/jM?�<A�]:�@!�-����m�k�KDK?���m�@_�'��;2$qG�]�D-�X&�ԏ�\F��i�h�F`�=��i��U�����z�2�q�����QCg���糄/�zd)�h��Ґp~�"q4S�G
��Q�t%T���ry�N(�Ǫ?�r�z�f\j?�'i��]�����$fi�e:�&0�~/���*����B���q��du�W���|���}`��,���Tj�!���{���3�9���Ë����+���7�n���WV�	W(V��@|o�6N��˓�\;
��{��uw�9����<��[8��si��e_�?O�y�)�q���^#������rr�#h�"}>�Y�� ���6���o��l}��Y��i�EM���
Z�v�G�h��恓��{ӥf?�-�/9(����5{�Hِ!j_�e%i���AC�����<���J�샛�d�1Z�t,E-�h�)����K ���M5������a4w��@��s��F{��ȾI5�C���G�2��܂xr�ŋ 
^�X&m�H�6a��#CGB7�(�f s�Z�9|^:�=��pH��F���B����7|�y�%����+�0�|�>c��d��7��~�B��d0����;{HsEQ2�h�C�������?��h���PލZ��ӣ �<#1�EǋI�r��Df�^� ���R��	�Je|x���rq�
��1t�6�Kp�X��'S*.W ��ҶX�O��۽&=�S���ƛEg�*OASA��u��N��9g��p���3�{+��_�
/�_(��N�Ȧ� ��,!ȅ�؏.L���X�lܳZ����Η�>�����QA_���A�U���W�Nq1�<����+���'TN�X)s.�M��m��<��; ��yEP�I���_t�#H�*�3Ӝ�{��lq�����P�<�����ppL.�Lq3��皥y��=��	��5��k'']���\��lR�����J7��}��sC�vw���-�&�(,�xR����K��=��-8ϱ��Π���Cߨ�H��#��4���K�T'1ZP�H��&KuX�k���;4:�<*��G���t<{�y>�|�J��eJŋ��R�7}thѶU8��j��6��*K�` E)�F
��,�K��P>�oI�"7�s>���]����w=�R��E�B�H��SO��x����᎛�������t�yҠ�݅&�C��*nMܜ�-�,���!v�c�uO�۱�i@��<�g�/"1��-��m|C��q��R����	�ҩ(/˰u ���Y��;w>�����������,��3�{0�@��[d2�!��B����m��v�sMD�]���g5�����j�jF"L6��l^���|@��!�.�w]t'�*���b�`��Q9�����B!���$��5��t�~�Ϻ���m�w�	KyUZߡ���ۚ�\��l[��#e�Zt�ű�J�i���g��Fj�Js�Z�ㅾ�B�-L(�����po����e��U��b0�� ��+��Q���D	�� d��_���>G�MP(��,���1�^�S!q�JQ����1���V���*��j9Cݴ�G��? g]=T0���D �k�S��S�}��G[j�v�	{��P,%��kϕ��Al6TN�Ci�*��D���~"Y�+�9�f�ɫP�����|�����a��6 �vMO:�5�V%����_?\dLJ����T��+N��<$ﹹsH>�Ѝ���zKLq��:�u��u�����
�\(�ӏ�?[��]L��@�{R�����S�h}��2(ߑ[��r`��zv%����>ўobPj�&�T2�I��Z�lh�T �f/��p@�N��O�`e����Z�8U?s��=���4��yb�-��|��s��k�1�"1���i�KL�?�' ��𯍭@��,�,ђHü����S�����,vK��:�ޢ�<�;)��v�I��0{�ق��*�مJ����X[Jx[�,�o0Sw�If����|���D~H�0e��ȼ2f��,�'�m�s����$�eB����}r��*��vk�	���FpS��ur��uv��[�YY
�#ۧG�L6�V�c#z\��E ���ϩT�!w��i$�1n���6�ժR�u+}�yC�A���۵^�E`Va�'��M���(��5�x�Z�׼�*
|�?}"л!�-:g͈�Cv�n�u�p���c� W<	����lr��p=fm"TCI!���*�ϴ��]��Q�l���ˉ���ey')�A��RF���n:�|]�t��̝� �|t~���,�{5 ��sY$�z7Tlgal���H��~�����|�C�evdL�j`�8ߧ>�<4���t3�!�#�z���?J���"�kH�l!Ҭ�s��2�S��LM������d���J#���F#���4ڦ6�P��*���رM<Ojc�|'����K�E�pٕ
���t>A|S��V�uA���%{��8^��u����%����h@`���Ѥ��zE�`-�t�0��% �t��]��+�qV��0]��	qv��6�Z�����\�I�O��~{�3
��\�P=�Jr�Pgo���mJ���T�Hb��7��^��p`Z��Ur��{�<�e ���1W�+A�գ&g�4��D4���(���Ľ*�����݋0�%D�$'��7�����jF�"'��kp{}xw��v��\��0}��vqTS�]���+�Nu�/?��.;���m��&����c�v�E�yO�~V��8�t����>ʔjl����u?ٴ^2R`�.��=��@+��D}���[v��n#��g5v���mg�.]G�Id�H�dv��3�J	xb(N :�1���Zr���F@y)n�����JZ�̸H��.�4�4����gA�͛�kD�\�����K��\��:�7/� �Fh*�+1{21��C���PYV��C=3���#
��L��2� ���E�N��E_8����r� \��¾
�ED�v¿��P�R���}(=�Ln�=7j/�ID���e`�ͼwj�F�%_5qS<�)G�Ƿ�{2��oPة�/Ҧ��Y��h�
�,/�pH[y���
̋�8#�Sp�+�p-ׁ��� �>�9�-n�X��b9�9i
`R7�e�L,)iXH^�)���+��K��O�A�]d�%�<��V{C�d�S���������*�g�SE�0�׶O?�j#)�p���DE��9j�|���G��.kB��x6�
Ԃ�J��� ��;��]�6�sŠ�`=���
uT��U�7a�nJ�W��Y_���%�g;�.����y\0���9y��=�����Zb���*�}�.��;n��c�rx0wYrw�7�U���TS'b��1�Djc��px��*�Ŧ�!�!p���t�^\s fK��,ؒk�ז��i?���L�>gLи���gFK��D|�k����)���"���Q�hJ��l�ҋ=�F��9Rt���("Y�T�V/�mzg��b��ɸ�����k��>��\��w�U"?���;�$���4]��	e��ٞwP�s?���������+C *��h�S5z��M�~��o����L���z@�F���,��^,�px��+W���f6s�LDu}��N.�X1z��u���εzO"��v�m�QevT�	.��Тmg	\��X>�@ �h�s�K��������͕���i�`0\�,w���{=�(�"�B�GZvO�N��첦��u\p|D���|VjLH����ޯY���)y��Y���r1
�\�e��+Ǧ���t����I �tR��ۂ�	�6�]a���%q��`]Ƣ7��[݌������gQ�>{8����N�6[@���(�M�����_/*ۖ��f&�d��K���<�xح�$�-ǛVm�lZ�W��B8,���:���\Dդրq�r�*w�ak�ކēܮ�-���!o�W-����N��A����TR�TM�'���׀Ӟ�%f�{�~V�m9�����"��l��%mB�S��*����(X)�[!�~�exuP0��s��ݡ\n����'`��)�:���d��ΰ\٫O P�]�������.Ykj>@�r@{���S��wW R<C_�v�1�?!91g(������?�`vA��좤���pۇ1Aꁌ��^��o���C��/
�d���D�}�+�@�3?���l���Y�6���<z={|].�<6㸫���k;{���Z��æ�O����|E��jO���+��7-��B. ��5�|�%��Qi�g��>)Dm��Ed�F� �t�)�X�y�W$Oa���Ǟ���"���G_�Y.���WH��ɥc��sg9
���˳�R_��9*�e�x*��t����C��=V0S�n
O���dS��\V�pMJ�* �Q��Qd�w������f�ݥҰc弅���� _p
I�`to�@���N��v�������K��I�3���a�$���f}�V)~p�G ��;P!c�о-z��W��@�'��I�q��5��W��=LGj�*��'`>|A�/�H��zD�tm��,���"7B��|=��K�y&b�����R�Cұ� �I���1H��lU���.��ńZs����Ҳ7E ��
Uޠ۩�/���liL�C/(�lS��p�#��a+���q��MV:�׆�|���B�!$x��wj���`O�d1�MD�����N1�ف��`�������K}�ѭ+m���eM<�m:~��V��i|RIH�*/.}�6/�hs�i'Whr�&�<Y�5y]8nV>�kM��i���})���QVM�G0�Z�
�X=�o���O�ng/]j(�d���d��U�
��K�K��M]�yy��=^p���ͣ�9����9l�<M��)�h�q��Oŋ�oՏ���J��;A�+�����wѵ�]���XI��T4�7q�E~�{`E�9�	X�w�ZOt������p9ĩ��!v	����8.�o��������&��v�?Y�c�*��9}L�ryN�b"�j3���Q(G��K�:ϒ�ft���ʔQ�0]��vv7�&MO��b�"����������|r}`�M�s���?�!��AEhC�b ]m/���y ��kJ=>�Ms��086�P�P�m���5��9��?���˭�Z���.���ƦR����AV�㔢�T�_�]�_���ew{���E�d��K=�\����j~8�da�S�=&-x��vUS
�P
jC�6%��4�Y�ݍN�&�5X��!49GH�h�@��ɞ�ncP�f��K�������3�+�>G��B�)n��E &=�C,��ӽ�O� N���V�S�s��lL�u��Iˡ����_
Ġ�g �+p���lm��)�<D|�1��7��C\y$�n4Ltw������,�������.��:f�0o�ۖ�\8�!��s�X�]��^�@��e�a�'�Q���҃�UrL<$�
�s"�Znv7��br�mV_�@�=='x���x�9
�^�
)�DD�ÿۼp���pGF<�i_O�ӔH� uV�s��fPƀ@F���Ώ���/h�e 	պ�ш�j��t�^�t�_&y�X'�qR�H�Y˂1�G��4~�&{�%G���X��j�a}c�w��}M"���VTґT��yN���9�q�^����G�����w|�I��')Iy��?;6o�U��	��F�U����r�kO��D��:�h��H1�� +!��> �\C@?'Ů>uG��Yep�ZH�%� �d�����A"Ͳ=�h�Hq�T�������b���^��c�߮��vh֩��ڿ���Tٹ�9�t uw��5���׼��)��L���QϾt�C�[PG�l���������M�֞xD\���*�xh�7�e�iI�cz1b��BB�ټ�H�J6�
Z�K�����_Cn������֒�4�=�����v�m�u3���Y�*|���q�?nT�Y\0FC����E \ob	��ؠn�h�ݵ29/[,�L��9��J�F�bM����5�VV��ZH>
~�u�����`6�춝�:l"��Ϲ��:7��D�vYy�=&F��ëb����JP��h�[*[�O�f�lRt�Ћ{�h�֞�x����z��M��j��y���nS>��A�f�/g���],���Scz񭜭@�P��MO�3�S9��������7r6{��y�hkf�����a�`�p^�K���~A|r��p ���h�e:���W��k@C�v�B�p�/���&=���y�M($-��8K̃���%A�C�]��������#(��Ğ���p�ah�{��8�䥐8ρ}�cE ��)������Qz�w�Cr0�F ��D�!���"��J�{F��nU_��cߏ�.��/�#���������}.$dU1��Lx��RTRj�;�H�FA�����s<oU�wjZ���a�Ϣ<*=2���
w��cLU��k+9�T�:�v;u����e4fe	?RO�\O,� �l�v��*�b�sŃ"WI��i�S�F��m��������]�Y���(�DƭZ�%N�S�,�ҳ�Ū�.e�YPMfޙp�c�9��1��|�w�<Ѽ�[$E+��V�/\�����͢߀��͛�ɐ��& ���XZh���k�GwV��)�U��]4b��X�~�7�~������Nj�1h��K�(\���Pd�~a�X��ap}7+l>�][4Qrn�CE�`�I�u��y1h��vɈ�VK"���6���!�m��!V��9�&�B�'�C�OCN��ScF���+w�ԸcOI�Hf�"�����k�]3�C���В-�y�; �&��k҄�mK���ߔ{��SP�"}���H�K�H����-r8 �����+ �\Ic��4�}�p�@ 	c����v|L�g�G��;�$���g�
o���e��] �dM�T����iM�y��6�
�z'd��������L��SK&\�z/k�KMXI)���5���2瓲�l��:�Ekō̩�����8;��%�!�+��YG0�hӈ_sF������^px������F � �q�.�PD�n,�p7����a񑌮�Ͽ�ф�����DV�OR����!�������� q�"�4��o,�?>��x��͍������.���a�֓�d�Deͻ�I� g�!���hJ@�������i�O�V�0�n�Z_�{�&��'���O`����w�
���D�ՓX��Wnr"�c�!��a䘚%P���_Q��;0�X�q9T�@�V�$�<_#����j!����k���ĻrLn#rs�TY}�)�+=��g��F��.�;b�_���ɔ����*�
E?cm�� �*a;0=��g���z�nQQf�����[�({3Vrǋo֛�C�<0���΁��q�l&e�k��n𿛭��i _���=�!���؍,��X��.��k��yev�p+�P��k�k�ag��ū*����z8 ]��X�0�
RLQ�kkk���+J'ԭ��	^��* c���s��}��[�W���D�D&�?�G7��Y�k�h���@��hB��,�>-^��Uͩ�ŐO�ގ��U:��Hs�gY!_�!ҍ�O�����No���6={<V���8 �ǭ��:��d?i�s�����H�Y-��D�A��nD>��P��	ָI(��6��W��~ѹi��C�fX4���	��d����h�c�qḹ)o׽o���$������t	j�BY�b���؎�	��A��A����_�,O��[Dd�H�v��y����ࠣ�E��;�0���¿8'F�p�1m:�ܪ�2�:�����NR7q�x��X;k�@�a�D�+9�\p���_U�Gfq$�����V��\c�]ZQ�@p�Ӹā�����N��Z=��w�E��ct��L����o�l�����N�7�!����������>� ������G"t�@y�3�oi��r�r]Ѡ�&;|�ߨ����*�"�0�=�ƅۮ��Y�=��"1�RQ?���P���xf�DEB)iq���2%b�7���4aF�r��>���^�̔�7U��g���j����>����r<��&O��Ii�;���\�8==]F�Fj�_o��ٙ �@d���ʿ��FdjlH���4�0����g���"����l�{���ǀ��i��B;Xj��H�����{��:���,��vXB�~O������t�r����h���l �\}�x�)���ǌB���rz p�24�aK�౴�2�x�"���P�/o�)1�֐4�d�I!���z�D�3I��(��v�{?�؝#=�9��V��tF�j�衋H9��1�����X�6�U�xy;�~�� Rf�A"2�o���h<���;��`[��s0{�����xK��/���h���Y�[0�<��6FK�-i����F�2�z�������5� �I�Q�k28�������SP'߯�ʂ��)���#���ׁ�iM���9�0n�i�MQb�f;��q�*����VǱ�������q�߯��mv�R[�A&�uca����A�F���^M=�}�7}A\�y��U�2�Ɋ��)�����D�Yٿ˅�	�d����v�--�~:����<5��:�ա����i��+p#�I4@�����kƚP�tԢ��ߏ���'y�b�^\t�dw,�s9)'�1��T6����e���s�L�p&�q�2	�$&z��fH:�TAV���AA�E�V��CIՁ����N0U>ڼ���s�xd#(Ѷ8��NN`�"����17�ٔa��WE�#Ǩ�@6���,��X����ɞ7�Ϣ}��Q�S����l�+�\I)}�4��`(�Cr�8�<��#��(=�V�m���k���@^������t�4c=:\p�B]{��� i�>��OņUWj��6פ�^ҍe�� ېb*f�G�]�n� Rqu���Q1����� ��r_hg����<��6�4c����N��3���ʉ��O��J�m���G=*����+����3�I���z=�,3�9��zO��.z����?�e�����u�_����t_g4r��C93��U{Z͗���˴GL��|6���Jm	�,��(Ś#�<�L��iQ�_��aBrE��}���jѠ�;`&� ƤV��0�",%c	���W�?q0&u�)��K������5B�bЇ."��+�p!� �M�M��Q�Ɩmw�M���}�s��kj�:`�5L�6����,a�r��8؇�j2���}���D���_]��l�"��#��B4^�b!�8Z������'пVL�Cm��D���0�~��	��\�6��I�g�k#��rom�	��o>� CV)7�'o��v�o����:SDi�\��i��zn�����x)���Դ�;���Ae	g�e����D%���c�m�ZJ�&���a�p_���ON?�<Բ��fS�ds��W-?���'ճ���x�'F��I$�˪�$@��J�BHȫ�~�OE�y�-��4�D�H���Eŗi�s�0l����$�������U]!���	�kQ]ܴt�3��$�����P<���M�E�x?�r>��l����p��i����ZI@n%�@�I�;g�:��ŏ�S����{�+|r��R����������	���[�j}�ŀBE|�kU����׌������B�UP?����'tg�͑��3�����{LV2��G��D��׋8~)��Zݽ�E���]46�����W�1+U�����*�q��'��A>��kV��AJ����J��YfN�|-��ܾ�����;BK��חS����'�m{ɤjf���|�ތ}T�ɿ�~c�m����E�Y.������RLB�D��9m��s&t�1BB�9�7�CHT5��SUZ�'�ڸ�C�6��p�."�G{���m/��(q�d��֞m��"s_-����2�O)�[Dih��ՙ0)�EL�6x��������P�w��!��2�Q�:�:U�>�!ph�!U����]�n��k��Z;���ۨ������@� �H(�P���ءs"�T�3��B���AA�mI�Dz� 1[U!V�5T���X96���'�'9O�e����/��`0)���S��u��5+jM��<�G�Ӑ�M�'U@��sZ�V�&�����@m�,?��Nm� ���rL��+�103���\w�f!��9��[F����|Hw|�v)1��q0�A���Ҝ�zpf��V���Q~.�X�.z��p�\U�_NR��L?�(���O}�G�Il*�B�s iC{3"(�"�]��H
]ҽ=oCђ�rFlW ����`�p�_uRw�����F~�U�ƨ~0�����գ4D�~&�]���)5��(��K�*yy�bs/#����vE�'�5d��D�^~t�AZ_�T ��Tc-J^b�?nk�i����U���)����'s�g�	#h����fQ�t��H ��H��/GSj��2h 	�j������2���7����KW��VkZ��;��'T:O�ɚ9\ȸ3Ms˵�����}@�H�I@x��U�G���U��2#��P����e΋�I=JN�A>���]T()5���[)�3��Kdbf���o��}�:�%i�O��=��'?��B�2�#��Ӄ�W|��_~�c��yP�p�1&�X;�=�,x��__:S,�t��&���w�P�'p&+k��:%�\f�L���+pw�HM�a|8#M��D/�:�^p�q ���!�)8;wre��	Z/�p��v�M�������h���K^H�ކ~�&ׅ�Tn��xr�I�B;;]u�s5��W��
�	�n�£�����g�}� �9���&f$��d�4�	��@�_.;��'�Ԉ$�9��=/��P2�&Qe8S�B���P"��x����{�ea���A���f�D�h�!{�W�Vzp��}Ʉ�{���l"	�#�pB���ïl��+��Wo��d[�\�ͨ���x�e��H��>����?d�R�O��$$��Es���3�뻵��3���gѠjx�F�k@��v(N���7,���۶�r�җ��^��G�%Sq٥GGF�į�\�����P�o?,Hh�C�͝��'y&�-����M��d�v#��6�ДŔ7ZT��Fn�e��͊w��~x���\�n�d/�#s�}h����_���f�n�Bh!u&*b�J��1g,f���F[�g,����bP}�O�g�\NI@�;3�P��W.����s+�]m5an0�N`���o'��%P��?2�Rޏ��2�<n�8Lֳ��E�I�_�i��w�����̀vm7����k"��s�s/6Ixv�{���/�Sv`i��o�+D�N>����0ܼ��
����7��Y62Q���D��\�K�"�c�,;�������m�$H߰��.�U6�_mJ�`�D<3�=�D���ۀ�Ͼf�-_�<�f��F��<�ֿ���.�F�͈�贽Û�Iӎ�o��b�J���sp�g�x"s��R�y3��"@�v9�!0]����#���w�4�wi�J.|�.�|���{H�`������<�T��	�ۜ.��#
�B�baR0OwW��>`P��t��^�.��==D{f$�(n�O�0�U��" ���{�!�>s���u�1����U���Yz�����F;�LV[��	�׀���}x.iXf��t̷W�^���yZ�3��2`�߯�+�!������4����J��F_V�!�@�i�{~_v��&'���P߬�e'�a��ԋzV9����"����e,$���&y9��l��p�!fZ
��*:��["W�j;BN�`��ف���V�����G)�����&��C}�(c��rۜg�t�����Y��pj?�Il�I~t��gѱg�D��H_��4��bF�l�o�W�zgW�[c��'۷|`p��^��+dx7|��D�XSs�R����p�m[�3�Ar���yY�h����9]h�E��{�O/@�2܊F��@"Pe���!\��fՙ�c�s%ӣ���j�!�=x��S]�DGt�p���L�����7:z�0n���T�U����xړ@Iܜm�9�|�jn�����{�>�7Ҍ�4V������yf���p]#)���)�)Si��Rg1��-���qNY�ߜ+Kh(�BFOU6�^���������W;��3��53�R�G�u�����Ŀ]~���,��=B"�q旚�6���;��i�5��rm3��JL���0M��Q�B�r�?�%!���ν碉��m�+.��:!u_���|�]�n�Z��֟��W�1���(��]�]���֊0'ە N|�N&��u�Z!˱��QX�7��T�o8E����2���n�UF�����v�±Ekc�\@pɄ�qK�K0f�,�b����	�g>�s-���1�(��{T�<_�ak���"F1��Ժj#R���jx�߱���8D��G҂�W�1�Hb����N�:`�Tr�f�k��8�z�f�Dx!-�E�W��3]�=4*6AqȘ^�J������x�W�wD�3��=�+��+�G�r��x9����o~�m���Z�=��=!	�b�&Ȫz����><�2���]\��t���˪���:+�E�!�*�O�YJ�
��(����Lm|e|�ԟ�����C������)����>� ��W�}��b6J&A�X�`&a���|�9�Ӭ|j��������<�`{����new��_�6�ƍ.oC�RW�ס�MaH� �_8(5��i���O&�(Uї�\Q(�a����4o�KMz������K"C	��G�tq>���\W0Č�����c:��q֤%lñ@*��A�9�Zn�܏���ZU�.R>�����}j�g�G8��>�2��2LJ�f �����zb!�QI�?�XOϾP'�5cC ��� ���R�ڨZ�k�k�gd��gwm���������ؓ_�^�h������&�G�A�EF4���nub#��g�1X7܄��?�7���H��o%[Ӹ�{9_��W�ssIȀt���Hh~+��;�T%5�d<�����o-e4�@Z�uRWqF$E��b�8.z^ <��j���߷��+yC��m)������[1I�]����ҍ�
��L�RY�he������ K
.�?|�~O����L�I ��-@�'�2���nUv�v3`n��F���r4؛�z��=�l��أM�V6�.r�R�E����l��A��A�~��D��<��@-f�v�IM�gK��	�X��d�$;̕�w��-P�+�3<���8$h�a嵁��<�T���������o��d�˸�>���w����D%��qv���/�8���ـq{��yI&����ٌ,{����>K�Y��J�M2�����%��P<�n������[��&��=��y�i�U������x�H�b
�^L�;`F-}�L��6� ��v�3��nW����Q(2��PdI�l�W�q��m^i��Qw8,�a�>A�N�7�ɮ}��0�1L}������Z8�ى_x?K@3�9*A&>�A�V��w��g��gh�y�D'&��/�%�{�)��T���dp*}VJ�c{j�(q�,*����Cn�=��@�g�
�ZB��u��UH��{cS΋&O�����ٛ��o��� c#����+h�B��&��C�o;�B�	�� ��I(+�a]��i#����ۙ��>;�Y�)��hߌY��'�K��l�f��p��e��_V�A��+O;1�y�����B2`�8�!@Mqh)��f�i#�uMb&1T��Wo.=�5?��<����is��䧳��/K�h�����=I���~v.m]U��	�o�a����6�j�� R��tr�UFQ1D�u(�ϣ!,������*�,wѴVAfӷ��o �Tc0_Pb�\��.�=�􏔬Cў�d�����oj'8&�5h1��"��;�~N*�tQh��[I�kWK����	�
����i~�	Sp�R:0[�e~�W�g����R��!����,�++���¦8-�h�.L����ʋɚ������y@��X�?�y"�w�L�D���V���@��.^j^�,�p/��#x��\M���7�nC"�Рt�SB�;��t É"TbZ��n��sٺ��_e&
s-O$�B''�m 7��_ݐV�:Zis1в����Vё���HoL|�s���<��x2�O8g��Piwt�#ن6�8;�KkM�h `�\P���U�e�Kx&����\��j8�):z�E�^r�O�if�"(2�a�����"�I�I�o�n=Ҳh��nu?i�!�e�;�����W���r�}�s~ � �����XW����F�*�$�%G%yE2��}�z� I�J��&`3Yu�W������:,��	��IZ�#>��Kؿb4<wi^ά70�K��sW�s��A�գ�I]��&�ٮ�S�k�EOT`v- ���V�M�_� C���=�VĒ�8C�\��MJQBg�v�7`Џ� `IQ���#��ِ�8h[g�4g�5WZ>O�?ū����,�F�)�%
�>�������a�WPR�*f�����ť*�e��C������Eƪ��/Q-*
�%fK\g�ЁS������ށ��ڹ�J��'��>{�r���Ajq"�6~��،d�_b��P^�p7�0�3����ȾިjbM�FA_!~���\���M\�`$E�j']���ʞ��?�,�����f�DF�M���N�H��C���G��5���0b��Q��	�~#h�����0�2���(��A��DO7-�38���k�yi4��K���cKD���@y'JE��#� g�XV,oSF46WD˛�q�¯�i0�	�J���F/}�&V�avЩ��Y��}/�$�� �����<{p8äQ��>�tv�SH'� ��+��8�<r��f�5s�X���KA(�y��(�֗/t	�d)����Xɽ��a7SXO��+M40F�2BT��c�B~a�^+:ݲI��.�CR'�'h�f�C���ltc��e�6�W��R(y���#Mԫ�!�?��j|�0+0:1��c[f=C ��=�t���M�$h�{���O�zl�(p82m6o8���몴��~�a��m�Syµ0��P�7��,�<� K�VVORq5��f�&9��G����� �k�[�CZJ��6 ����"��6CA��3�:���%+�U�,���ʘ�����X�j�y�?'���׈��O�-�:S_ib���_H��~�'DVT�;�e3O���X�>���?��Ij]��oO!X�'�pa���ԣBA���e � k'Ù�	��A�������+�ҡ>�����i���M�0����e��*��t�Zga�n�~Y?�5��L��3��_���!�QB)_��Ɣ�E�fa��\C��	��;�To���Ǥ���M��[��ր����GA'�WM
��_��4��<�6@=O���D o�O����`��.%h8K�'P�&�Za�_qx-�#y����� ��ZQL�b�ބ��R\�伾�>Bn�duae�:qc�H4�4��b������'nl��^n-?�s�;��9�^e�P �Ԟ�m���aK�Dl,c��y�/�������pqj1�ޕ�%<��Qxcq�(�;)��J�l�̂����%T�b��+�@R��ۚV�B���UK�뺁,��!����.5BԊ��!�U-�K�����PEs0V�ap����'}�-"̉lL��z\x��2��@1��keM~��l���OB�u�)���qыо��:�4=z}��x�뽞I�k��+���D����m��\�s��L���is4�\�*�R����j����v^�:(��6J�_%p��T�5�>T��;�ܫe�'���j$�ٓ81P�g��mlEd?�+��?�������ꘗ(֧� �
w�@c�et��^������$H����ib<d[OY�62Ia)��S#zU��9��u�1U����?�9Z��̞<���Th0�|/������K2�P�[ Y�.;��3j��ڔ����X�8�����x���"WIf���1]W�8�h�Ū�1.���J���E�����A. L,���۹�G�K�n�og!��| �,����/8脓�����HDXGAi�vx=�"�7.2��7�]qc ��d Ϩ�� �J��?��
(i_�@�F�{1t�62�j���w��]/1e�k�k��%����L�`�7�#����@�:(�\�&�4�~y���� ���Ό����g��"v�'�����}A
U;���OҴ}SvMR��������\�@�ş2���Z������`R���E��#{�<��s��W1�&��l
k��?����MA&�I)�佝j�Թ�<�>}�9�-/����K��s�?ZR����v�����"U��H�GA�	�.N&y�aO�ٜh�)�q��j�L��5�o�<�똰 �N(��Q,�3����.��ܥ�O��L�O��3�$�W�����R�a(<G���JW��0�1���#�Oh�p;P<����W���dx� �}��Z��Gx��@�3(��$ی��S'����9�黝z�69�	C�@ԑ�\������XhC�^s_��!��\��р������2���\��ܧ��!jj�B�F�o�U�� %��3Y�X=s�:���Q!�H�����0��RΎ�"�n&�m 5b��:�j�_Jʹ��<��A��<��6��P�^�]�S�h,�Qj5r���h9~��)zAm��z�>4>�:��YRp6�,#8� ��R�H�u�7`U*F!d��[XP�I�/W;�-rY��|���me�b�Q/,JiT� kM���ږ��W���Z+Z�vV���G���~�fFvR"�v�DN���7�9�xH�g����b}�������j�{�]�ȼj�7z:w��1Y-��v8�����;V 3X�/{B�����p �2.A��-l�f�,=<�|���At��ݏ"���T\͢,�:%n���xN�e�8R�j�Z°�#�U<u���$p���>�
�a����X�j�w%��zk��7�y�߼�T�R~�/Y�R�!��2���'�5c?�#*��=E&�D�JϡQ0�C)��8S��[es��^�,�2.���n�<��7	�m�p�=�v�ց#�y�>�w��ݻT��w�wk��S3���.�����P*%�3��x�6[�)a�]^#���㻡�=*�u�|I�p���y:��E�^Hj�j��w�\�HŸ�]_�.��!���~T�R<����da�~ih��mb�\%�Q:M݊�ٖE�c�)˃۪�Wb/��!�W��� %�N��2.:�OUor�ZAXSh@��$S�@��re(��W��	�F���
@Z�((�V�O��!v
[sk^�u�/���Fa��ê���?�����F�|VHL����ߡ
�͕O�C$J�>3ꌐ�`F{��7��ci�&L�^g��7&�� �˫v?����}z��:PU��:�ϛF)�S��	��d��&��{>zIO"S��qHFh�f��7�P�u��gm%s����x���ϝU�������c��0sb�����G��h1UɎ�A*&��� ��Mt�8S����lk;�]l�q�w7h�� 8Kn����-ZU�X4��F 8��F���� *�	��<��������2�/���M���c�n~1�ٶ)��GO����F@���IS���8='P�A	D̞#�s|��N�F�m&��8%��]�{Ռ.%��W�qd�R��d0Zp��	[Vg��!�|����ݎ�Bn�^z������1�$�h�WCvm}8�1/���D�/	o��=�(�r�e
���>�����n*�*�T���?k�OM����H�P���q��q!��׽lO^t���M�TԔ<.t��=R�feg ��;-$7L�I�(qЭPɍ蓴����c6����������#�.�zb_=u�d���"��z�>R NF^��y�8��^���U@��PP��%r�q��(�
�T��3��W�~5����D�(�Y�{�
�}�h��W����'�-{Kls��n��U�`
�J�'t�7I���7�Z�>�_��T�DV,��^kÙ����e�L��"���xEwSZ4iaW�!�Դ4?>�P��VP��2������q9|�)�z�"���O��4#g)\$�}���ԭ��a<RT�3�cr�S'��E\�ZG�7;��K,�3��$c��
x�B�0��?�|̡�ͦ�"@�Zo�(� �>���=�.d�>{周�_�l۟N �W����5����M��(O���,�r*t*�ՙ
�+�	�J���y{��/���!%t�e=���:=�mQ�q��Jn\:��^0��5k;�Wq�Јv��i�^�|6��K���?'�d��A�qV���� }�Q\)I�߹�)[�
�v[X�Uvm�?��X��ǒl�J׫�(�
�(���n����]�.z=��1��t�P[[䥂��Ji)�8�p�;�<L�v�p5�Q��5�p���r�lP�"�KqtW� n���w�vy��Izo-��#z��U5�:tt�a�$3)�RfK'?�I�Q�o���������@]�bn=�r�-�V����(5�F�����吉 s*�N�I�y�� ��h��V��l�	�^��b�*
�ă7͉���ͯV4���ˠIz���p7��|BfCV�T3}r����q�a��@]ʑ9;!h�\zʤ���<����U�oH�a�,��{�抃y�$�����-w�w��^Z[!Y.��wA�1'е8��K���ܝ�s�����۩]'l���տs�Ӷ+�	� 6da̗,��:v���T*��Jd8H��(a�;0xf��jϰ�}Q��d^��B�0A���C��_���:ϵ?c��u��1z��FW�u�F���,N�cUR����[�"4�n0��<���;C/�/�Ѿ���D� 6��{�q!k�Lz|�o�ZJ��Bנ+?���!C�1����tG�1�l�(�Q�B��ՙx�hӀ��t���9N��WU��bS>�����O�o���O�4i7����<c����D�0�b�؄����ƜK-BG�EV=�� �����]�����_E�t<�:�Z=�`dڝ�'5Nn����sB�Xa#��d6�B|lZB)���K�~ǟ�x��d��#uZC��(V�ri)��)����[֙Q�A�o�i$|�b�?���Q�2�}ĢOai��aE�V��쮯<�@B����0�aeq��]_AD4,��V�R��.�'D������pr����OB?�Mf���b��7�z�{~�ZF�c~����1AQ�g���g�FxXN7�	�D���`��(�>��M,E����S{�xP5�֔���e-���rhd>����/��W�Z��>����N8_
`R$�n�cU�4�}���2�3:Xv�y�k� ��͕�뉱t�;++{�Qo		>�+�18�n�d��6�t�����t���RD�SkI�un3y�!��b˟��e�#?�y��pu�=x���EnHkP�~}هw�Sr����ݫ��������g.�g�&"ɽl���� �a�\4=nL63P��#��>�,;l34\a��MQl��B3,$*����(�	 ��XMi��Fp@8HۙH�~�7���~�����V����0��W�<l��MZ9YD�8�%R�5P��203v�/ c�o�p�{��-�<*��:�~���L�_�9t'�{�ꡨ�A6ӫ�9[!���B����‍�̤u�"�K�Uz	ؓ������>��� �J/��.GZ��=04|�v/�͙��"�%�5�r�|�>)ǉ�HC��$`�H��XBo,�%��T��+K%��C��1�P�P�:��}O~�^�E�t-܋�o�%a���ɽ�)�X��Z���ǑY��mO��3nNw��9甥~�h��!��d�ק��UW&�B�yFn%W@����
�)8�&�}�9L��-Z��z�^���5V֍8w��{�r�Z�g���t!f��r�6�~TɎG�z�A�tF}�<�5yu�e���U�f��U�2H:��0�\ޕ����n��]�c�1��u���i{ɷ<��I!_c�߆��ko�G�kL�^���\��|/N��0.�]z�T1|�p���U���M�������5��-ʪ�,��bS�)+Z?�5�h	�o�i{rA��B��s�����i�1
S����qL�ף�*���Ͳ�{�,E3��c8�� �����t�ΐ�1g|�p6�����R�n#hߛ ���ƫ�yp��U�w�X��=$T1�_x��huCq1��7�yN��L���[��[�^S�Mru�ɶ���Y�J��|v�U�������`�Ә����ߢD�6L�4՗��
�'�P�*I��RqJ���t�%= �BT��Β?���@^���;��yM�}�^�� Vs)�wC�&^t���#��ق����t���z���5)d3A���cPʔ�6����]K���Y'Av������(�@���h)�
\Ӹ�!@����w��׳��s{��I`x�Z���E�'�F��PD�FZ�'%�4�<�� 9�"f��M_�1C���=���!#�n�T�젪½۵px����	�X(p?�V^�׀�j�	k�g�F�a��3z��� ��P��j�����>����$�|Ajݮ�����c�EΡ'1�$�>b�K�������|��6d�"f�����h���A MH�k7gu�$�fܮ���#�aǕ����び��m��7Ӫ��N�?FQ�oZ�W�k�`SW�8f�!,�_�ZC�>j��8��֨��r���}�[b���衭tm���K�C�Z;[���s�������*^2����wH�2}:��Y�SX̞��ޡn����+��D=j�u����~Z��h������b�����Z=�n�Ys�O/SD��  /qt���B��Bxw�$Ί�ǿ*#g�P}�+�����#ynB��U�(��D�Y0�����ĔGuB�M�� J��Ҩb�>tk����^����)�pC�K� ����un7z�.�Q|�r&����B�kp��]k/Q�󻞓�S~����U�HD���VO�=:u?%6!���e�ΆJ��/��,:�"�ۗ2E��0��Gޥ��o��=�tl�{�N��f��+�KE�еzwQ�<�s�&A+�4j�Mm����K�A��7��1�[�����3��&z����7h������IB{"�m\��w5�A���cry ����HZU��na #>�� ���u�	 �ҥ�ރ�[��S�䆿��g	�蜷��ה��}�G�p��
��u�!Y-n��e�}��V�̷��)*��&zu�]g�< ���.��4�L6��4<Ģ:y)� �c]�6�d��wC%�^�n���i�VB��"m��T.�
M���o?(����5V)�[���;�=�IM��N���]�J�����4���s�mB`���1�H m͡�-��_�t-ݡF�u��Zb���e�j�i���(�ޝYZΎ��>�C]�k�w�X�$ �`��aS�y��$p_h��蘝n�-wU�yx����׳1�w��1?��/H�Aۍ��]�O�ްȬ
��`�[�����룆G���G�s���b��c�;p��yמ���69[=��i��J7�K^fbܞTb�>f+ݞj�p6���[al���Խ�T��FeS���f�'���g �\|�C�B��u[�ԋc��A��fF/�/ o�do6��*c���k�	�����ti�=�����]������A�`��'Bneb�e�c`dp!X�����yc����3R��:���nI�����c�C�њ�ĺ�u�!!��v]kB!�J���A��o�X�	�ޜ�@�*�A��Zj��DɘKշ��	�]�y4���EF=C� �u�V=��'܌�]w]􃕇~'��Ӓ���V���~�
�%n�t��t�J�+]���Oq�sbi�����lv�H�˖�߄Xk�/�(�����v{�� G��h3J�f�F��zJ���2��2Tn(:p����o�2/���c���B\�EԲ�w�x��B���6�D��[�}�<<�mKD����71��H�7?�%:�yLSF����K�;Ͳ���F�Q��<�RF�g��Ӥ�����\�9���:Fw�H��ڀ�B69�с\�#�ł\!Ÿ��7dNhL�I�.�Wn�y.�[�;�~��A�^ԅ~�A�Nk��Yd��(<(�������:w�D�!:��Q#��~�cH wNލ!�.��6/XO����T�Jw�e�@و8㌤K��p��W� ����m�����LOx ��hI�_M�k#����������^���DV;ȁ��>3<6�	(؟KB[xÐQAx�3��t����¥K�d�X�g���.��^CI@5��Y�=����kY=���}�=lCM ]���ށ2��Ƶ�6jZ_O�p܇�ݏ�*��?��"K���j�q��I�⛳u���Q����y��M�Z!"8��]'v ^�=�s���|u��+���HNB�6�BwD�qk3���i-��m� [���B��ނ�eӧ��	>c�&�k���l�劋t� �/���?����R�CF�6k)jWU�r�c����F]}�WY��^��!C8��h��n��`��������U���j��%M�:{���������c���LI���#%k�v����*�l/����n�~z�9j�)D�)�a�[��b;j"����ˬ��U[}�qS��}m���u��H⪲ށ��%����i�K4zx�k.[Mg{�����'`�kA��x����D,�"�|�2#�(m��`�Z�%P����~�YA�pZ�~o��8���fdiZ�W�>M�����g�!2�R�{Wy�6Nj����6�8o��dw��%��6j5����fF��
G�G<H�:dˇ&�u{����`E��hi|7�������@y�S��0���{L?W�q�;Om���p)\"���o撣�t� \ʄ@��B�\0S�N���P�4�����x��}-4�iI��f��%?C�q����7�©���E=���%�/��z9�	׳�E		aC�� Ӊ�{C��8��ܫ�E��Q�b����^3>�J0*���e*Ȏ����@@t�?u 3�G�Š�~W���G|�� %h|���R ��tF�f�v�y����1gO9Fb�?j&�+����Ӎ�UZ8���c��J�;.̴����
@���y�4��r_~�(���..Y�E�����}ރ"D�8���U�Hϝ���76��t����es�&�'��z�
��"_B)��X�B��W�08:?U#X5�����u�|4e�!�}�>�y��D`��(R���S�r
,�D��+W<A�P�s���)��n%�.�+Ms��7§Q"\R�ͳ�O�(�¿��g=��Ɔ/�b�#3�]|ݐR�
����l�|{d�nt��2˟�bɽ���2Q����I��!��g�4�N�${�m�v����q���s��(�r��?:���Ö�{
?���l��I���� B}7�@<UU��P�X����]y��1��k���H7w���e��]�˶iZDB���I��Nz�\U�Y�H*��H�����W'���[uJH����y�|�SjH n�ek鴋��n�^�����:�c��^��Jj��L�6d.�a�UL9t���	��)*������̰�x����uL�k�	8�[�oYq*�h�˞�c�n�F��w�P�@��$��w���"�R��H��;�zf0�
2��MgN!��K7���'�vA�n��䖲-�B�����)!�V>A��I����G�y�5P��k�mT���IMEMkh��$�I�p�۳��9���b���4�
���KU@��v��J�c�s��(5l��V��<="�#��?��]5�`�l�s];��
	}��!�/�C �y������B��34�#R��~g�%�*g!�3�˴?0�%�/'�Y��/>�Rey�a����K��J��x�\��!\�������
K]C[[�#�#�$a�Y�KCY����/��^e#Py����n�a����EV �SP0�aON��1�~��X\��i��%�M�|ͯ�鶻fT�fR��rT���w�d����`�p79^h��P��e����	J�F�uֲu�Kq��9�8j�џl^���K�����!*g[�Iӧ�r�(k߸���,Du����*M1�����#�	WiM���8f��P����j��}sP�k ����Xc,�*���^���AN��+\4�wi�L�Z��.!Ɍ�0Y}L��EY�E+����M
8��ϗ�z
Z���'?Yv]d��^�P��H	E�gr��Ư�,�D	��XT~��9�V�@|��{ֲٹH�ΐ�����+�A��}�)f}&x�@��k���!-�K�֑)wp#ǩ���[�^�U�+�+˥0Lc1�1�c��y�~�^��[
_V�>kX�7z���yx��V}B-Qi��O	�M���! Z%m1�O:�����7!Lfl8��:�D�T��!Z�������R	Iy��!I9ʙ�� �8����aHa�����\&�<u�a�`��"����K+��[��.�Eji���8�̊�����K
1NM�꣚�oD��9qͰU�@���e�8��r�.�#��P�����"��nމT����c����tZ�@./��]��}X,KU� {����Siѭ~x�re��D��P�&
��K:W��4'�q#��b��O]X�v��+��d=m��=��rǢ�,���xeT1�mK����VC�������+#�|5�����Q�[�\������1�zI_!�)��}����u��/�
�A'�*6_���l�kʾy�ƫS��\�����p�����}wl��[�Srq�[��q�����~�Z�L��E�jzΔG��ջ����>v�c�R���1�?ٚ���U�4���ϸ�4�K�5�J9�r�{Đ�$L$g�=��V��Χ�;��&~j�g�6RE��q�˜A2px�H��#���L���Oz�BjmӔ�Y#�펈���~�xp�1���8����7�*!����SK���tbQ�j�w�� s|�T�+�/�²�"rf��Y��+%��hk�����.�*v$Eqj��.��,���`l�^�X� ����;H[�u�sPReݚ�!��4�eC@��ȋ^Y�z���ٓ�
�๷�C���n�[�G���M�8kmJS��.L�V�;Q^���&jy�H7ȧF�K��W�⿢G*2 y�u�\�1YVq�iD,�H]��%N���
�#���ϙz>q|�w`�Q,/��Tb�Y9  J����.���qvu��DV�#�pW(�3���/�x�*��=sj��q�ݼ�L�P�x:�.�<����	mAo�Ɨ���ځjD��{"Z��&�`R�4�(��X|Y�R$���^ �}��W7�Z_Fx#Q���u@Y�q�U���2�_؛}�f|)��K;�,�>Kk�u�⯙�h����+��{Zƭ�z!��ZE����)�Ah�paK�)��̇����KŃ*Y���6�D(��.��/�lEG��n��G����d*4��b�Zqq� ���oڬY!����a&�*�e�]���y���1I{��C#C�v�2&_:rIoD�i�a!�$/s;�j���4�,�T��"0��[5���������C/�*읜>"��tq�%��:�48�s#J�9:���NOыW>�X�u�v{#���eA~�wZQY	=s& �����-�=Yިw�;�5GB���H���t#/�#�rt{�`�}�g�1�Qo<�>X��p͖�#d.0�w��GyФ���(�#�9�>E��I���#�KW"7<8�nA�n�R����1L<A���x�:�D�n�>m���_&`ߺ2~���h	aN���G�xHKmi��W���J�@�k�o�H������m�kt��/�'�E��Y�Lآ���l �aP���oبU�X
��w�ȑ�����N-\�"1[��;��IG����fU�q$�Pcgh��9I���Hǋ���8h[H��'�t��M�����v]x!����b�͑�e�F���D<�Bj���\k��fd�2���_hQ�RV~_�m8��6�FJM��	�@69�T6b[�c���e��s��>I*�r叩���$qJ��bݢ��2P�.��eTey�h)5��<��0�Q��9��cӰ������X�{����F��:f.j+����Օhk��*D�rӖ��ļ��GDzm��JU�z��{�bC�����p.�p^�o
�!���m�D�+�Fڭ���3=�^WP��R�ak)����l�8��9 ��v0��i�UrG�R� �(@s/����#�| ��ف�2��N�D�n�\s�����"b��BW8ʥ�b{Wq�ȟ�P�{���;�N�O��G���^}��pдa^�c̳���5v����M���%F<)�Lf{4�0��r�|!g����d턨�߁��i�)��9色d�k1�5c@}_v@�1�P���* %9�"T�����	V�?��ܫ��jb���l�UG�V�XR���yz�C��T�;���ȟT��h��CM��q�x���RZ��e�9O�Ygye���h��>M���w�SzĈ�K5[�%}XM:����Y}ɥ�gƼ�t�S�ӎpk�2��s��A�*�̈X�R<Nv2��n���B[��p-#�o[��nAs<譲>Q�G�E89�����2p��c�hʋ���
�h�k�)���|�U.֮��g�I+e�b(ڒ���sƌÕ�u��Wc��s:(n\ܖS�ݗ�;�D�k�L�*,�a9�D�ʛrO%�O��K7�N�E۳�*�U�x�c9��6��3@�q����R�Z^�+��r�m���%ш}��T>yTHv/r�"՜��ʵ�1��8&�'���$��X�4Ka�H�\�G������wS�񕨤qZ��v����P���~;�FQ����`��Af��8J'��&���WN�ːr��@\�Ph�d D&�0OK ��e�;ǟS{�:4�� �3eF|��Q�M�[ �r�T���}d��7CAc<���V׉�ܮٻz}X��ف�}%�'#�W�!$z/@q�O�j{G!��n�fs����2��
��P�o�*�|V��z{^�B)/�(��[�-X����Z��o3̌tm���~�3�'&r$�Yw���СvA��l��$�2E���e�@��e��pu��ۣ��O�\�Bz˖�[��!�#�>��KK�}�����x!���Bbx�;�������!��jҮ���;�%�?��:�~oy���ɟ%�1�#�����@^r����=g�q���_���!�c�I�x�n��`I��Ȗ�Օ!�H��D�pV����]%�$�γ>ݩ(.h����Q�	3V��f����������`P/b=�G�R��D����.�]5%��&J�%P���8�g�����[dPE��#���k� k毿UѪ6��,����]�!�g�,[���&O��^:Bv��5���txI3V̡O�m׹ �ȰՖku���fF�+=�߾�q�r�$�ReV�����Y�/ϝ�D�N�o�]��a���
L�hP���LE�><��zѭ%�6{�)�^��wQ؊r��07�K:?3L���6¿E�y��&���#_�(Q�[Yv��\"Ě\>��)J���i~���턕'��A[���=?��􈏡p"8���~�X��>�v�9xgN3���yy+��l'Ⱥ�V�������vB%А�2���"�e�$�V��P�|��5���q��>�;��*<?�xRq,�Ԝ/Q#�w�ч�_>�8ط �%���s|�]?�Cv�A��c�����7z�<������f0z���Ƀ��5�֗�U�/���ԍ��]L�Q������qV����2	��H��uI�$j�]�9|����c� 3ڱ���7�$�O7T�]�o͚м��J3e�~W��u%�q��d�	������8���iQi���ym�5G�#�����{�f~�@I+M�	���ם�ND����]��^��|������[�$�ڏ�)g&轜A5p��fwApT���?��P�TX�R�t��M�P��&����� �G�$�90�j�{��Fr��4��ޏ��Q�FtA�F�̀����F�au�E�'j�Ϻ:�ne��w3�3,˪a��Ȅ�\��ϲ���&�А���H}Ǳx@7�*�h���AB��ԇ(�R�i��2i��[�Q'��3<�&C5� ���EA��kk�2 +w:��c�\�-�&�]�s��yt��d��.E&Yx��
�R����*�6F^K�ݴ���0���!��m����T.�[T=�p.EHUl�Y����u���j,�	���k����7�?�߈�9�y��&���8��xy9��R�B�-yf���i_��L����Ό9;�����K������Г!�W��.�Z�R��$��H�0����/���JmAL싅���C#�l$:U�͛���[ݵ�n��֟7���F@�p^�_�A<5C���~��-2�؂yZA�k�$���2V�d���Ʒ�%i�%�}:����u��+�H_��$� �ä���J��gd{O@��_������2E%�%��أ�6�)��a��ǎ�����}���D^[b��!n^����:��@��9PO�(�Aˈ	/����!-�v�*q4?ؽ��ܪ�.f��_T��w�Z��^��N��FW��([ϯ�a�k��F[�<f2O�������8q�щ�֢Ρ�jI���M�a�փT���*��7m�v��iΘr�9����p :~�I��	f�t�x&Q2�ө}��ZX$���e�Fg̻1H��9�[�7�(T�3I\�#��:�r�oi���U;�����&g���q��ymM�Ŷ��T$.NV����3.�	��E�n����ӈ>A�Ҫ8��Ԉ�亃g|�����=A�s�ob��/j8����$��!�'�H!�,\?R�Y/1�R�J0����|p1���w
���p�-'�7�����Q^���Q#�Ԭ������-ut�>w^H5�����h���������<�[������O��m���۽h� [�bB�g	�s��5ߟ��#3	g߶�ĞN-���ϔ%����iCWZ����I�`U�Q��1����G&�j��_�C˽���s�;eW��x�ͯ�^+َ�rM�ý�����+���	�_��%��>f�����'�a���7�ґ��#�S�Q�^��I�3xI%�W�pP�\�~-�>ϖ"`�BF�鏎����>�^K�`˱w���Q:9[�6��߁'(��e���h��?J3x�6oun"X,���ԝ{�*��C:o�,�y#�K�2R�+���><_D<�������{�o&�����ex�5���P:\�+u_�˻�~��.�>u��8x��>p�]i���-�lt�>�?���CI���r�P=��;�i3G�gV�nD�S	�{�h�*̧-�iք'�8V����N�h���| nmi�	������[׃nMД�aP¼V+�(hz��,7�Y'4K�g�{_(eT���O�zNU�����$�"ţ�h��~�DD���� l#������:n�V`wUu��X��~�dϘ��]�#R��$/�I���%V��?R�''�;�S�=3��5	w������v{&� 2�T�91���w{�v,h�l�؁	�bΞ7|=i�(����J$�{g�V�rG��27��w
���l�9����6nd�n<�Nl����|�j���J��W}֬5�`k��k6a��L��E'�k���
�ⱘ��4�I5���� JuX`F�ϲ#r��ܾc�E���<�@yA��D�f���^�j�<"G@ˊ�<���m�%�gɺb����v*t�w�8ݵo��!�
I�a�t�Z�6��[�b̸�w�tv�KR,�C�Q�y4�J�iۀ�+�`�N9�Q���q�>@�b�����6����[���c~L71T4ƽ�"ej�
6���1�ۀ�S��	�u��ޕ߬j� �cC���w���x]�B#7P?�	*����C(mx��$S!��v�D��:U^^��p����T�;߰��
:SV�FN"/��ό6V��jiMq"fyyY�vE�t#��Z1Չ�1V�)/�����lo��P��	|y��rp��j�)�1�����?�|^Ҽ����AWGJ ��a�J�h�pY��VS��ӝ ��\ʨ�N���3B�lj��v�h��T}�Œ���-�3 Ӗ>�����w����S��ӆ����W��NG����В�K�f���7��J��c
��^%�Vi�
I.�N�4���y���U"\���L����A�a�o���?�|z�"2�O�^c�-f	�i~u�֊J�����K����$W�q@���p�1V���w��-)���R=�
���/�co�����\�_������OO�]��Yt�jX����}Uæ��T(^F�WK2T��n��B����Q�t��]�3p^��t�c;[��jL]�]D�E�>z"w�����fYH�E�Kpm�]@�v��;M\��}�P�΂�g���.�U�'O��r^�{�iC h8�t�(�Ӫ���#�dp|R��O|.��m����ҥX���V�Q?��F����	.z�cn��"e�ٙO�R3*\���{���T��6�6W�́��=�[��[{�yi���N�/p��.�P_�	�aP�ln��w�w "����Mk�2��e�d�|�5��@Mn�����\��13^bgp���l@+`i�ƞ��@�Vm�1�<� ;�8�'�+G�a��`�M���#�l��-���ux�R͸L|q^`����|�]yo�h"�c����������X���B"����R;&��wTc8��mm�p�b#��I������tq{�wNo�U��0�0g��
��7P��ƄP
��D!v���̡V�i��W�^�;bsv�S�?�Q�4Ǫ�w͈%+%�_j̙��\����U92�.Y)yٔ�����	���\@fr>S�O�l��[8و2M
��'y� ,���D+��/$��ƛ �8)*xw�2��$�Ļ0�4�/�p9���?�6p%���C(�C�"?C�4�Ͻq��n���'��HN�&r��ђ����A$��Yptg-���uB� t�`�0�]
�P��&�g�$�4Muu���e,iq�ìJר���H�h�B�72"��@GFf�t`ʙq���Ov���C�]�}��RN^;���^�_=y�c��x��}�*v����tc����Ť��	��&z�x�Y/�9����m�8;_L�gu��|��d-�j?��f$�MO�¯��w�T�Lƣ'�^��b�n�3*[��p+;^g�]З�`���3�YC�ĝ�8����AD���* ��/�~%��j��J�����DԷV%[~����u|f�Q]�l{�x�X��W����<B�"��2��1���A�:��&ӡKCMO'����B�� //��N�u��f!,��a��!g�$j�ajUM�<�� �8�Ė� �@����n�ЯjH� UQJ{bZ�} )#�-_]*�x�,�; ��t�θ4x��э8�ɰ��������nY�^0? /
eh��
7�����l�Q�?��U��W�J+�����0��rr���w�\�S1(z�銺��t,�}E���8�j����D��mE�$�9֋	�"P�4�r��8JU��x��7���E�-n�*~��v�]x%�0���(\�3mo�V��Dr\�l ��Zɸ��ζ��a���):�Y��2�f	ԳJ�L��(D�����;<Y\�ه��;�etA�+��n��t�X��!�6#�46��c^
�*���&f�LEX}�_*�27������R4�	�G8Ϛ�fH.{�'#F�ū�b�z�,l
�@rl:o��[�|��􏋲�FH�ڣ��ܓ��F��Ƞݰ p�ֿ�b`X�Da��<L�[�2�-�;@�d`<C�Cͨ��-�x儋ӑ��%��h�vV͑�o��� X���� d�ʋ���q��l!�W17*����?r0xf���!a��S4%�K�O$B�����˽v����3��aj}�ϰ;���������n��}���r�[�N]�d@I_�ܤ�iLC_�b�v��)��2�]�j$�/ߍ���̏x��_�X'��J�@�|���N��<"��ֳT'*}x�I�.f�w3�������x�Q,GPP����G��q�:��C��g�������&���Jsqb{��z���V�X]�����Vja�����o 5#{{��}�_�ٶdGZ	`|��i�p�Xu��>ex���X�9�W�+᧖퐌#\ӂ�q>�'��/�~S��<�Ζǃm
�ڔ4��~5b��i0G����~G��$s�&��<�����L�V:��!����aK�4�1%�} ��w(��͙}����b��o����Oٚ��ڱ��Ol2�`���.��WW��	�0��t>+���Y�Z�}h�b��N��t�ah�h���Xߪ_+ȗ���g�Z��^ {�Ȫ��g��H��C�3��q<�<���DS
����4*�$�d�[�M{:e�=��Y
*�N�#�,��.!T��(9?՜cv�n���|'*J��/x �����fws�[��W,�	�Dq��+'J����8:\��	��ջ��M��ϛ�.�Dc���q�����e��(2�S�	 �{�G��P=]�q��8f�u���� �L0��֓�e�f{�c9��,�Q�5�Ya�s�T���4J5yÓ@�G�i�9�y���c��Q�Xfk���5�>��X�M�0�J�ȷ(�Ew��h��8D*���<6�;6Px�wa/��lE�"�$gK�	-3P���R�;��İ#���3Ȭ�йw_�͡�/h�L'�m�,��FΦ�H���X�Ց���չ�h�]�.��i�4c���F��{��u�����ޮ��p�Yt���Z=�V`/������1��O�^*�u
.
�|���Rƕ%�òU���0�@k~���;�Pru��
���A��a]6"�"6ET]��O��?�E��Å����N���{�o(e#r�Q@��^��\󯦮lE �kZK�$�6�eU���;9�6V5E\0�B�dB)�;��G�rH�M���Ñ�9?�y��E�\jQD�fU�0I\�͔���І�but�.�Ž(z?0�1�"���2Md�-�0�!iVm��u�L�c�t�E*;�2aY�Y[cz0[���p)��4����tՃ�d/ר.=e�p$0�x^�=p/t-� b	��9�%���wJ᠞Z��]�}�T�`G�h��$�&5a=�æ������M߂����%J��{����>R��)��J�N59ޝ�evȽ��ׇm����MQ��k�̩�D����E`�-��r���W�S<�m�|#��ڌn�C��[���G��䷈��|qv�o��y�pT�LEH��b�?<kH�l��DW4W�T�M�\�3�CR���*�X �^���C���?��<���4j�f��s,$|c1����i8���l#/�xj��\%6�*g�r=ʧ&�}x���7X=��Fl��I]��z��]t�sIg��b&���-9���YC�N�o5R9�gZ�3��M�������8����Wfn�Sٙw�O	Wý���c���Of��'u�h�q��lH����p=(��s�;cf���Ok�<&�N!����g�Ĵy{�\�k@P����Q����;����=��������z�A%�p��(����g�A��f��L>�+6���Qu�i�u��u��	u�;ی�[L��*I���l�89.v���)��h�r+�R*�vV���ˑ�sy���i���9��%L��y��/��[������)�y��`<�o��I+ȎF�׻���彔{e�Y��������5kW�@��M?r�.��U���G�����lDx�����l��_�2(eh�|�9�D����S��&�4]�V�9�'�U	�8��ix|ӓ�9�?��b�}�'j0�\?Ϳ���+��.���$�Q#H�6���6�JN���]���`ty+LcfR����,��­wՑ�����������ٮ뎿���՚����av2@2�8���`�3��z{�(+��*�?�1��F�(F�|�1���l��"�T��[\I�T�+��b�W�G�%������
�&�"惸����8�u�h�n���˞Ҋ"?f���s�y�����e��5q��o������h��6JE-�_��YN��2Ua���;R�F%[�v�th�r��>[1��� �z�Yf���'LGif���H�!/����m���7{7��o��(7��C[!�=����d�e��تۓ�	3��
�뱋�=�Xz��:��� �6�o�	9X'� �l���D�3)&�Ø�:M�x�
O߯���4Wj��&&?���kԱ�Z�G#�T
?0��;1čP�;��R'�I�2 &TwW=�)��Yw����9�풪	�6��a�]G�����?'����(S���O��*����[���[�~2x��v4��7HnZ�
���[ȇ������M�Ŭ2�.;��F�IK��\(_���v�+ݟO5�1����څF~��.�F��5H���$5�T�|>,=��
I��^t�9�L^ �M���*�V��FՄ)����1��!J��!6�	Cxn�L��h�	:g��#jz}a��{�$���c�:|�Ես��c������<C"�Y�>�Kk�������������t῕����7P��8��m�&-���@�����윻�t\�8�5-�����=��h� �����p⠼�d�����Bw =����F�h{ ���/fɣs�""�N��3�4�����!�����S��jO���Ƚ�`>B�~n�b:*z��K��� d���fh5��u[�����#xj�,	3<;Z^�w���#_�o����`�B	�@ym�O�%���[�����U����%p�
���;���Y�(EO}KN�V�F$�#�,5�JVZc��`ى1s�z�͇D���C6N�j���KXr��,��ŝ�L�������R볠��t�4Lx�2��ŵBŞS�b=�<b՚�Y F�ȡ:�U�����p��xڠD�t�ko5~?�kj�����D�o1.�G���wZ	C�I�O 'z��xOc���X���0���g�Bqt�|L�p���r_n��~�|!s���2�$_0�������ss����F�IG)H�^�W��M?�v� �&b�� ��$u�s�y)p �?%.�i��u9R�/�\��紿�\�C�>�I��ҷ�`/ʻ0�:O��NN!�~{��!$�^���g�p(�ax�׊��<��Tz�e$?DV�3�$@��oA�OK�����ZW��t�a�Q��������4���=b�Ո(��
�ͅ�N���i]0G�$Wx�e�	h8�Ԑ�"�
�{�"���V�U�Y8hQ������:B��e�X��\#ӳ�Q��27�n�?f��H��.�9�>,~�>����䦐�*Zw�����l4]S-Fb�2kE�xYX����6�-g����,��Z�/3���hm����D�A!6��BAC�S��;X}�`a�
iG�)ƾ�řl��H/q��C�ʿ�S�h=c^��yeIE�z�1g�/�.���۱��D[���彬JǓ�z���>Hs+6�Ό�'J"� �~<m�r����N�g�k����ln�/�#]��{N8��6�Ԭ���*�s��%�R��#}[�x��F��N��I�r�u]��rn��U,Ȫ˘��:�3�h���G1V#�f�
 Q��G7���k+�=���Ƃ���;���1�DŕS&��ҨgƜ�>GN�DF`dY��.a��V� m:�:oU�9��Uǳ,
)7�1|TI�~��C��F�4�6��-\k{�ڨ'JZ�H9���<����0J�-)���)���΁<u��BD�����0IT���mvԐe��t���C�'���F�K�F�������g4��ӛ.Ǳ�Ĩ��O�����X�|�B��6g�=��W��Y�4��|*�S}Ƥ[�=_��;-O���>��'��}�`��h�ق�8��S��<�)jNO�"s�w��S/�����v�L�������vL�[�
��˶V\/	��9���Z[8�r	�J��	�пc%��Ol"?b��N}v�\��i+�H�k���qQ%'�E�Y�u��4�fx��$X�@](<U�Z��߭�_K���^;:e�ӂ0�<k�M3�k77i������AY���FXf]�B�\ZH�I��T��	,�:`-՗�������������(���J�CM�]K\���qY���E�>a������X��=6�%�x�a�1H�~���5�*sr�D���u4�HSɐ5�F����L�1b5�	��ibn9�d�!He�o#��>�����(L?7ƈޔ3.UXY���tZ@���s�U��kۄ��4���WD3"~�2�󖞜%��i�?���[�5)g{�����LϿ����J)�=���N�2����a�N;䚤�1�>����ma�8����(�á���f��w��@|]�h/l�?ls9���r��A��\�u�@���R���<�A�R�_˷��%��B-[l���٧��ʂ��C�j5��@ ,�O�e���r%�&��������r���$
��������w\��ĈN�'�=���/���dɾ�h���!��#��څ��ʬl��-�	���y���O��^�],{�5]:<J�	��}�Q�k��i�uX���D�B�n��Pzc����C��,��Z��E�zB<0#zk�Ѣ�E���I[�J, �=3g4����LWN�˽Rt;)�	�	|8�ej���b��l���q�$@�u�����%$����6��x�Z��:d�	TT���9'��*�ҨP�Iw�ᒿ&.6S�u~'G�� �,U!� �����A�u�iL�t��K�&cl���]Z�F~Z�#���!���k��&e���u����t)��Hɦ8�������N[���1ԍ5�j#WR���s��{�v�>�|�X_q�Doxu�%O#oȿy+D���a��vW���M+�=��*5�j6�}�?*Z���7��I%���E,U1Ӹ�ɥJ�Tk��v��LCNx���,��(�T��p=Dw��[��To����W
��Ӄ�J�t ]�nb
>���EM�S�Z������kl���P1Є���;Ph��'�CB���O�X R�ȶ��lZ�9��D+��q��Wg�z���Ժ:�f�t�v5"A��r���m$X�c#�hҙ�ݭvTG$;qd��4��Y���2f' �_h�X�K(\:� ��ԫ��@c�L.)�WF�7�sg#Gk���IA�86ղO��>e�U�UMJ���������X�Ĉh ��/�m[TI�4�Nlׇ�xh�M��t�N�({�>���������:t2_d��J�EC�4ʄWr��i"u&P��ƛ�ՠ^`���k��#����0�C��
�(Caf��, 4ߞ����h��<�r'v�{h��MZ�#k�jXXSx�ܢL͊9J/̍_ a����3~�* h�J�C8U�cM�'6�.V6߫^�|�Gq�h�X~���nMn�������88��[Ncܡ�o�ߒ���;�F��Ԛ@a�G&)%���Y`Md��M�`��0�T��2��u���P��gX[� �x?P���Um)��k�H��r��4��`��Ti���)�6�����|���>;��U����g���9�l����z"���)��+�C�rK�n�-`�R�M]�<���h��u)\'�
|�(R��O���0�<�d�fwV�{=��Yj^5�_[�UA3�mr7�V%Q�f�L��Cy�50M8����=py��dj��Mk��n
f��Hܨ�$��u�ڴ��%u����v�Ͱ�xI����h��ů�{�����螩ٳ���_:���Ȣ�by"8��s�!�/ڂ&��*�xx��qz��aA@�X?<N��c!F�EH���nϡ�O��d���htp4���p�oF9r�˃�-�#�=,��ӓ�I�Hj	��1�����p�Fs��>�6��#�����g(�=�}u�g�pY���K͇��A��lς~Y�����;!m�БTT�P��j�s�W �*�r�����X�,����AN�Z���c^���,:���D�E�
�Qd� m���B�z�[��rHU�]�w>��(M��(��8�T�(%Z[V6��'�B�5J�}��9f�C&OS��[#��a&legn�_IR_�q^|M>�l��iQ��`��^�X��z��}�O��j\�"h8�G��5��#��9u~�LF��é_y~l1�/?l����@5Ef]�O$�����r&9��R���@;g�`e4���P�REg�TD8L����o�:�%P�M䡆#O3^P6�-��f�) ��O�="%�Յ�ӯ���υz+a�R�
B�t��s�r�L��*(H�}�����b`�����_Ȃ����(�l�j�5ۗ��DڬH�jN��$�%��	�"i@v���Y��Z:3'��7�b��1$�)�^� �nL�7�.-U_j�M��~0L�9���~:4������� L�]�筪ز�հ
��
��W��,�P�.M��>�XE�4�=�E��W�J0��ob�bzB�ŷ8�O�K�x��H��2a�*#�c6Z=�++jy|�?:�EV���j�Q_��ŗRD��z>�iF��ݿ���9fu�%�{��K2�b����1 �d!�2���&��v��HD��'�y�jd��o�=�JH
,}`��� �J��X�;�*ޛ�.,:�ݻb��lLN�̯S���Q�v"�*.��y-�>[��Y<E����P��xno����M_��a4�Z����=���x.����k�����U�ʸy�;�{�m^ነ�ξ� M9%.��Dܦ_>��GQ���������^¸ȷÀ�h�@�}ݬz���H�N -�l�Y�J�0��[�#.f�0��Y�hw,��j.~�0am6JN�as�z7F�.h� q���F�D�Y�%e�����eH��Ro���m�(#�<�������d�I8j�h�tV)���3��J7�U:;'��=����p�Gm�����W!��
���2%��M�O�]���E�Ю�%���X�D��-��jh���,�e���J����ϟ�����J|M*���-.*7��`�EAp��� 9�A=N��_�fH�����t-t��`��^D�j%������2v�ݏQ�	�����md���f�;.�];z��|��!=C1�(FY�i��'|�0_�?NNꄝt��U-U}�ƍސRݠ$��Q�r�,b�˒F$��&�[g���2���6AD@�iC��@i�1�+7�J�s��dǝ[��i8B�%Vۉ����h�W=�&�.y<B+e�r�1�{�j�h:}�B{�;�����+Jk����oOd��LF����K��v�1�o)g�ڜYi'�������z?��*�$�ꌙ�g'�'a#�N�����f14j���D��H�ѮW_��H2�x�-�]nv�&���t��j�]�^2�p�D����B�����t0���Q�2��H0*�@�dLU��nǏ�tg��A"N�H��$3��AY�p/OQ���,ե�}q��@yj�$���28c�,�O�t&-ܞ�b��K�'��.?
�>M���ⓢ��'���~���C��_�&�T��6�yi��5xg#m%�������� $8��;ˇR�P���X'�C�V����������oO�ݝ[D�`U�)�~����Y$?,�
^�a���amt����&���ە����kt��P�T@���oC�gR̊���05@F�[0^?2��=Q�~� �>�z��`���`Ekt!���i(7o:<0	�&�գ��A�$�Pm��x�������+�F�rmj��ex�&�5Ʋ$����[F��_j��	�	�B�`�m��)�<�	K�򁨖k]Lx�,�K��Lw�u���%P?$�U9lP�)���-XɈ�se�	v��ȹ%���#r��:P���fTL��}���Z�9�ݰ%�/�*�����g�QJ��e�$��\�
�刎�G���#g��1�x�q_�c�ܞ��n�V�AzHt{x4<z2Yʹ����L�� ��J==��^��!ף�q�C:����f����D���*�c� �滖K���
��:�5��0aq�kd���oNρ�Q�ݤj-���r����t�>����;>�gJ��$]�Ry^&��n��w%I��!S��9���'�i�o��|�$x��~��ȸ`��s19	Q���TJ��6�n_��'^���������+ݖ����H�6�;�$ �w�1���!���<�Մ���|�Mlۓ���s!��&�0�_M��<OYk�r+�QOG��~�:�m/c��"	k:�&��Ke%S�袙�q��̝'}��=��
|}{�ٕ�!��x�/�d���sᏥ�T&�Y[R��~����On���.!���]��!����|f�ڿu���+��ۊX�{VS�FQ�����lSPB�l�C���y�JW>m��J}��Ĳ��W��'���g��I�^����k��C%�����`�J�J��12�A�J��BB8��� s²��3��U�ydV��Mlr�?�|��4x	��'��s�8[ڃ�#����OeiQ(���C�l��x�q�-���b�j{�5'=�ҢM��(Ȩ���vn��@���8{x�}�x���=V�b4%L%D48���e�z*�pm��^QD:��r縀07�FH�ٛ�Ȥ�>�}�4�&����'����-��4đ�ܞ��x�n�� �j'`�E1 ,G��?�Q������v(p�?�ǎ
����<H�+
2������Ω��}�}٪¾����@� * ��z7�R�1.�>Ļ��;�$3/D�_ �(h��f9�p.+��#vk�`���Ƀ�ד��4��Xq?f-��'i5�sq;%�qc��з4Q������}���m���/��u��8ʆ]�!�t����T&���+�j8e|�x~uR@� +�(uw;�c���rߎh�+����|�? ��;�5z$j{��e�$���y܍���Y{I�f_�25�������e�*e)��-Q�/�aF�Er��*��e�ށ��x��g]N�0=�,}�H���6��#{�'o��i��s��)��V�Ḥ��	g~�U�;6��.V��%�%�ѷV��&j�eu���[���B�ήB�vv�J?�QG\^j8	gOuξ@�����S���=K��+�T�-Rӕ;�F[%H&=�{C3��2�W����V` i%Ј�����,���1>�w��bݯ����P�6w��A��Wk�;�v'�^�!�wI��&We��a�_!	��E�ѓ-���e����h�ȭ�F���O	 ��.k��-Z*p��ԓv�Fl~qr�YP�p�[�B�⸻���S�G��{��$�<����,��扮�,D-�*5%��,\�d���K{�Tdv���X�>!���<Û��a���� ��Co	���V���q"�rkb)������a,p�g�a,��WPnÏg�/�k��A9t��t�G��2����,P�/��_zۀ]
�f��}Tf���r(^6�N�u���aT�0RTa_J6N�ɽb9�Lz���E,�A;��n�5$�r�]7��pth�؛l�ȼ� ��;���U����(���"�!�p�h};x��qAjAT�q,޴��W�J�Y�������K���d�N=\�/1�f8P��x����&���������u�q3���?��?{�5k��V��@�9uk�^�bL˷=��)������k~%��2=Qw_*����:�����͊��40V&c�:`e��M��ֈ��;���6�_d��\�T$�a���R���n淚E���5<P���Dͮ�DDJ5�(c|Md��]���ֲ�>6�y���{�U��{�������J-W" V�|��B�4M�������E�b��b{W�X+[�ѩj���n�+����(�W[�b�*j2�j���pYM�|�j�g} lR͎*������h�[���� �g��eF�K�ӻ�!��i7�4Ś#X�_�?ji�f��H�� �WS4�7�Q�_�@]��?S%f����S慉lgi��P��A�At��h=Ó �;��X(���`�Kt�~H��È�t��~�?w�e�D3Nv��*�M������z�����H���X�n�ln���9���J��C��2 Q�	�V#u�|VPA5�!�	B5�Q\�'���i��lݎ�F��m��4ez_�t���f:&a8R�����f�]�����6)e_V;͒��3�?`�l�0Rf$�phA>V�HX�E0+��x�P�]"�Q@Ȍ�s�����X�9�gv�cf� H�}e8?z�|��*�{b�a�΋���]�\Oa����BW���5؇���g>J+��`_���SC�$UK�V��*�6ɖ���[׭#���*��$�,�:�@$�7	X�$4V阏z�}���H�\͏�L�F��:�{�LN�� ����6	�!�[���4"� ����l���;����v�e�9��'�D���O� 1��F4&ڲ=�6��睜�+�WK��$?�g�0~M���+Ƕ<����K"�k�āCȃ_7���r2BM��l��o��og��W�ЇE	��h�u<�k��ݺ:�P\���%'�Qӧ�K��K�4����#����b��>�78�R�wI�2�E~ّ6hGyĆ'$X�69u%'�s�md%w�]�OC!���DٔM�_'�����z�QA��`�$�j{6�̣��x����|P[���3����+��#A���&R D�"�++�ε���<�����)\y"�9�t�٣$��s�K��JD�|�Y�C~�׈$��駸W$8�,97:%��r�q��2�Rя2=�0Sf����E���[$�F�0��K�EO�T�y3�8�T2��l�w{R���^�1�(�Jm��9��o�"84kp�N���&�G`�M<��-gj�(V�-��U
/�ĉ��챺��u�߉%Z1�jI"�0^�rt�8���*��]r�kV�(�C� (��AN��0A���K����:}� F�Y��|�� �Q��]ps�����<^Bs�� D�<�(w OёD�Q�T	���dј;k�}�TB:�`����g���>�������o�X\fRt�`<�� ���>��3!���A>r3 ��`�yW:��-x��Z
nI�3��_+[��8Ъ��?�"��"ؖc�O������y,뺁�Q>F��tɄ.WM��&D������z����T	A�GD�r�1�/�[�qZQ�b~���<J�Qc�%�"�ax�V`��E���uU��2�k��Jh�NXCWe��Vh�I�ڨ�B��Gܔ���J���U��0�S�4ʟ�2��q3��*#�q062�-�j_�����<R��B�&�F�D�J3�ٷ$�y�;�](B	A�9`E��������u2�]����G����V0�A�d�:�k�A�m�y_���T��O患� ����O�k;$�н5#I/����dƕ#��^l�6����Խ���v��tAe�ǀ����+¹�� >�_^��C&�R��
���R�2v�g#����=U������$g[������Ig+���xp�,�k�=�"8[�A爞�T��zN������jD
�N��&f?LJ��X{g�	���+���F�.���~#�_H|гU���Ăf4<R�+�P����m�5m���5Kt�^�>r2��]���������\7�'��'��C��r�{��~�칚���������)�(���Z	X�pyT����P�5�?SQs���횅��a���J�D�$�T�,���ZI)>�#5K�^-j.�Σ:��/��p��cy�N܀��|&ď̋TЏ���1  Sxs��!RD��^ʺ��9�sG�t�3��r��}���Y����v?f(ї���	���i�P�Ht8��'�dN�(!�i��^.8\�Ø�%A-2���B+�}�F��윣	���Y�w��n�B2�6�(�F�H��oVFk�[xl�"
M��K�[X�(tHӹ���5uƜ�i��"p�m�#P<�t[^�N�c������P)X��*�Ī��j��7B$QK\�Y��A��q��5�Rj��j�	��9�?�B�	��P�Wu8�0nՍYY�ҾM�W��(B��*��<�`��+n29%�F�]��oa�E!�.a�E|\ʶ�\���7���v���3�eu��gki?���{�p���fN�0��T�bɲD{��Wi[���-qC\�h#V;B��4�Dh���7������+e=��;Z����rM�q1Li�S����0 ����\�z�Hė��7���9GMr1���f�\?/�Y����JKP�o�\�z";,��B�]��y	$U*������B�"y]���'�����c�r+&���l��l(m�٠�;�>N�Y�����^��F#3W�>ff��z>3OA����5��q�dT	R��>�G���\?���Kh�y0h�����;�09p��g�<�xg��2���d1��=��D�����~�a�
K��s�_=����Iɳz?~vn���W��[?���_�	n^�~��&S�p���V��L��8DJ��&"o?fP{�R���1ηL��@	륀o>[�Ãg]'�9���ȰBݳ�dS�dZ��M?���^���v��l�k�C��7c����7	�e>63z�G��>ž�;���X2W�T�;�����V'W޸�n�wZc�E���Q��ؐ�~T&��M:�n��|iB3y|Qs�|�zN��������H
�m���I.nE���5����:1B�!A������������(6ʋ@n}޻�O�a�w4�A;��E1o�� B/rKr��ε�_u�T,E�]��#��D,������vՌ�Z|�NL\\��7$�O-�\��,2�h3�)��>}wڦ�
����)w����Y� lb�V��j��i[��0"�b_�-���dn5�}�SPb�{a׏O�z���;j�s!V�j�)D�z �7I󾈈�9!-��w4���s�����jJײ]g ��GrX�!Pn�k30c���/^�j˔(t�PN�3ۗ^;�57ݶ���pi �K�0Kq�+l2Q}YNT� 	��%F)�t��S�9�#�I,��>�~��h��	QW�Ǽ��Q�L|+"��M�P��8�n�iտ�ˇ�	<�Ĳc�I�*ٵ��
c+<?��<��A�^�BD��49o�h�R��g�N�H(�E��[�L׮YG�<��C��M*_���n��r�x�)�����x��R9#R�]�L��Y���7�N��lzH�2�\�$_����9�1�F��i����ai�@�>9x�'�������ٽ�t=\��D��q�t��[;�,�]g5eY�P�s[ gt��n��]����,'B��Tbw�t� �?Wn�zw�od��S9Q��@�ȓ8d[	N��r��3�he\Tѐs�]���m�� nN�m6��H�+X��ʋ׏3m*m��G�j�@����:�� ="H�Q�����,�=�iV<�a
�XVU��1�`�c3籤�}�+H��~�J���	t7�?.�����6�#�<I ��ѭ5X��D��<�S+1h�P��6��yL�>*1q�������I���3=���LЈђ�(�^�5Ni^g��uʹpR^�L����+I=A�It�jd�c��Pm֡V0�<kr�P+x#��t�͕�A�RB���T_��-j�AQ���W�04TrF}t�X)�.�K�
�����|.V���"W_�SwK ������m�6�x�o���6�V�1�z�oU�MVn��x�z�6��AWU8G�t�����k�����Vg2��e�h�:��&��ߩ���B+gB�7�f�-�$[ag�yk׈�uK��!MU\_���ԮkOh����Xܖ.�[�mTX�;�� �0?��}�����H,������'�uF�A4zp����"��8HMj���Ъ��
d�/>�xZf����/�Kt��u9Ď�� �
�ǖ�e�����\�	��m�R�ϲp��O�n_��.o�ύ�O������n�0L��V�q�Evc�8���/�l����O9��s��u_IWJՐ������$'k�|���tӬe�E��E��ؽ��䦕i�-%>}�r�\��_�x��cEkw�~uػ�@f�G��b9gp3�!� �Y��qLNϷC����r�+�e��|ף��n���"�(h����C�ٓՍ+j�Z��:7ž|�J�L+�1}�l��I৏7��z&��[�(�3�4C#M4��?{�:E�9��ypxu2Φ�EB��U�ec����n��X="�06b���*���|�@\���0�I����� �@ �4u0W�F�u���[�=��2	�����l�v*Yo͋������|M@�d�v�+���e�O���"��F[gq�k������N�G-kp����^mT��4]S�(�g���+i��6���߅�y�J��3�C�-�Z�I��������X���^S^�V̙��WK����J~*ʭ*An>"30z�*�O�̒�:`����Z=����ݰ\´)Pw_2�B㍗N��>v����	3C��N�F��?(3q�=wt�,��b�H¼��$k��n�ha5CЈ�k\�{�����oQ'�ZH)i'��mm��+ �5Z2���BԌ0͗c3�1�����
#[@�Z�L��v��٨i��]� �4]�{�E'6�@���m���O �x�ʎT����2��;���Jn�6��Ա�¨`L&�����x�L?&��}��J1]����hf�%&����𲎼 0d/����D�3+���O�J,��=U�ߵq������{ެ��Y(�5@��{��ܽ|��|_��͊�R�H!m�3�
r�פ�t~&�7�Li� ���m��H�'˨�D�E �������fJ~^���5�'J�"�ru`��F�b�LG3�ʠҴ�Td��U�r�+ހ}Ӣw��8A�r�D�����!X����_6�-��_p7AY��ˀ��v��Y
j�f�9�e�;fX���$2܍9hp���M��u��0jT�B	�Ϝ�~ot7�AE/�BQ����$�K���#��E�qF��%�8�`�k
Zf��l,=?�_�q�<�}�5��+��#�fQ�<*H��;���.HҸ0���|��*c�63��\6߉�����\Ia�!w|9j���r��L���?�wK)/��`rV����A]ʤ�I���/<	��v�Ss"��1�nMAF4��&�L�"ٸ+I]���ᨕ�Wl}s�uZH��G�p����p�IFͷ����~��Rס�s�؉���{�6ę�*eS�T��0ztU)OqS�2J�
e�x���<����\���x.([l��'�����a^�>�;IIN��Ŀd��o�O�U�H� E���M��l��OnC�~����J���_���2<��c>�~�[������a���:䫬�x~�����m��	�ˁq���B�c�A��g���ưx��EX�����$�sӊ��W6gl�1�qÝ����/���h#�{���i��Z�Ȼ�� �"J��FA'�ހ򏎈�Վx�;��.)��֍�,�g�*v1|�C� i�E󠊺�ٻ,\�˼x!)�!En4�s�f
�P��2->6���*�B&\{[��0#L2Ů�Oݡy=�ؼ�#�VH�.���0�c�چ�x�nI{?C���~�Y��Ҽ�����
f�����)@7�RV�?M9U˚�F�DtY9��u�G�%�� M�Y�P��e ��AZ��mȨ�
o�z���j�W��9�E,J)M-qs�f�/��hoSJ8�B�\�or_2	��jb�$��B�׺�3ďPw�\d���-H�����91�H���D
�e ��"H��g�1�[$2���������{Ѳ6L�PaW����t�ЮY!��hK>��Y���r�#�����y�!��\=��`ݵ?h|i��v/��	����=k|�(F�وoN�B��˺O�s��<�R��ZB!��j<�5���*�OO�R���m�����N�Y��_�ɱ�N����(�ݕ��I��-/?	(N	ꕽK�!�t�o��~���ޒ��Ӈ�3x:"���Xg1I�#K3©ĩ�����r���` ����I��Uї�H�k/ ��$��)6����CYS]����P��R�T��ގ��8Na<�ĀKl&8��׃�6/~�����N�ŝ��#��%6��+O;���ˎ�������B�'�cp����N�}ll7\��?*ߟ���H�V��O.�"�]�����i�+�s��k� ͠��=>i{!lp���Z�9'��s�5����c��tf8T���}J�6����"��u����y�`���ewQҿ����#t�J㾵��9���d�R����H6}P��p>I������n�>�&�}�?+#�&D�&%��J��|%�kH�!�.�3?FL_hI�Gk���HM�A:gc�Nҙx��<a�5�t�����ab��WK!%Ө�J���W�ܮ���9HT8�Up%���lA
�Q=Ԏ����д�tT��38��n�4`L%�nW��J�4x����P�${�!-�w�v	:\f�ߛ։t[��5�F��'F��@�b&�O>]Bw� �peP#��(T���jy�d���\���5*]T�/x�P�3e1 �+�+AY�P�aVLQ�M�A\ 9h����[
`�@���'+g쯩D�7y����6P_��p�����hR�zr�;9L�+�mfgڄ�[t�ݿ�7�l��e��y_�M�������c���}�0"����������>�^ǋ^�h�u�/L�y��w���8�l����a�S��X�0dp���!��W[0�zM��m�R8c�����f���t`w�'̇ sgH�;�)���&=��"������j��Q��'1��W��hw�����V��5� ُ�S���ɕ
^5�yp3�L����wΰ��$���Х�#���BF� )2}�,���*��m�a'S�۪�����2�ύme�Pq��y�~6���23����=�hy��R��q�r��_x�.հo�B�G���aU�����}�g2�ph�� [-�ݛ:�ng�BV	�?�h�:o�a6!Nc�Lg�6:�����u #�1� !��랍���D�Hs�#�HCg��w��ru�����0���g�4ʅ�9r�5�;���1@�kw�cE�i��x��/\k�
����[@�(�8.�80�G�m>~��h��gQf|�� ���/�� dH�ೳ����NO�籭|]�E��̌�ŉ �u�m2I�Vl��oÇX��������Ƴ���r�������S���|!k�:�Fx?i��.���������o>
(��6���\�\Tf�5�f�
s�r�eG`��V+ȭ�瓦���Ij�HyA4��"ݞt$��M����Obf��nY�x������s��N������N`�m.&���c�2�ť������ڹYC���eR�u��xq@���Z���:�Sq��,�UV��^2J_MY/!���u��&ֿ���mͬ�aJ����0��/�?�R��3
�~�U�Ɠ٪�&�o}%��HТ4H쥶� 	"��|H�߇n�ݻ�SD���<?�Y��*����z��;�͉��UA ����C��(x�H1!�
z�`}	��W��W�����!m�M�,V��(S��@���c�%\[b��X���SF���%����KO�k=|�5���+���?Uu�O��
� XU+~��DLmzz��!\)L����yˠ�����_H�k>�� I�额p����Tx޽��:4�1{��$ {���FS�f>7Sr7{�Y�!�1g�sGZ����W0ݓ]�V�)����Չ��r�&p�$P�61��
9퍶��GA�+���RnK�гn�t�E0@
���~H�h�_�����<ž�A�LR��.�)�2�u�aqh�.�P��-Z�{�#�q�֢��
�����ܔ=�	_䩟*#�e�r<����u\H7=<CDݘ�b��`����#�r���{<��w��N[���5c4Rd�y�0��"�s"di�AlV���G5D��J#H ������eLj4e��.��ŭ
���3�E�l�"��e�́{��c�����6	?����X!�"G#����%C_�js��4~t���N�0�������9r���e��Ck	���U�(A=��
B�rU� 2�la�U��� �l�7.]cT�sٵK�.�(M���Ĥ1�Cl�l��"�����'U��`��I���;�M���<�Rr�����_f�Q=C���/.2����Pp�{��2�����⿂� �>�כ�J~���O��
���|��I�0���\�!Iߧ�ܾإT��9��/�AO�U�h��9�(&Cn��>l)��lP��n3��ݾ���*�<E1�����h��Aƪ(�nC7�V�ڣ�CD2�n���W��8�8q�����rb�hnֳ3�,�����㮒��)��`�����O�CUM"E�>�5�6���c�d�#U�d�ݩM]W�[@���Z���l��]�_�Js��\����ƪ�v��!���J!�^h��s��]�#�i�΃�V݆3]�.[���t�NC��i�h�l$Pix(�V���tb�A��=a�$03��d���C��ܝ/qg F³�<�K�|K�e��R��]��z���`�}{z�q�:܅���X��&�vl����X���Mg����}�#&y����q��0�6�ø��H����V��wߴ8B��06�k9���,>{t��L]�❒��Tgғ����l��Ȣ˄p)﷾��Ö���������<2-W=�a��%�DNh1T��I�'=������Ĕ��^x�0,%}����.��VM�"'�O����n� �$�Our�?���{
�x)�'��S��i'{�OK�����wI�@x����t�͏��H�Z�(�t���4���H}��k��3��{+�eْ���n|�I�4���?�{w�\"@y�c�c�P�}{��x����Kд�RO�Eb��"�����a�$"�,Ө��ZZ<2�u�8%O:��PenTE���o�̙��0�����>*�z���t������:��T4)uw��h���p�TS����V&�Ds;z��(�ʅ����O�qB+� �ޢ��t���_�����wJ��
�����}�.w�/�1ڵ�{g0�wf�>f���_3��>�l��!?S��4�����������ZHS����W �:�W�s��1ŕG��N�'������;bQ�����9�IY�~�k�K)����XK%�t��c���;�q�k������S�5}�y��#@��<�ﲫcX�F$��u,[��6P���Ӗ3���	
j����-a�6�W��w]���,� �O�/g
ꟊ�<7���C���2�{
^�ߍ��uz/���R��4�>�=!K��v��>&���g)��X�},*�:]���K�r��I*������,r���GȲdiC`�8c��g����44�aU�+Gk�����8��ᗭ��d�ׅ]~Y7����)Pg쁃��@�m�u7��xU���D2�_���[�f?��d�;Qߓ�J�X_��nٰ��}��	�,�G5v���T��P�ה�ۿ�ض��?�Źڭv#��vN���N!j�]�����\��݆�`c�t�[���d��y������x�^ǀ�'�ے�\NV*�d��Y0�uO�t*���q�b��҆��t+�
�?�&7WY-Ŵ���fb܊(5V&�7	7�����R#�am��V�A����>���5�ԟ��nH��J �y��sw_����� >}g��JmҤ��h�߲��q�go�Z/��8n'˰�[�p;i�����z��������K,��E�* x`��7�Eޝf[<\v�i�Ob�	���j�i�r���A9v]ϙM�2��fe�}_�G�'H���e|7
�$/5B�)z�у�˻Ez�D"acY�5����M<QKߕ���c�դ=I?t4�����4���{T�pm�;�Qjq���S����gW1����pod�.���)������L��ŶK�ٯ"�w�,"����/-C��vL�@�'9��=q��ڦ)�oUM��C�RȐ��p:z����i�g��`�Q�r�=�����4�Jۜ8F_��/�	���ܤ��t1�i�Gf�R�+�.B*���1�a�1�p���8ֽ�YQ��6������J�)
Q��c�8�9��:e�V�a�M�Q��3z�i�X�it&M a+W�a"��ڬ��Y��8�	J��S�P�E���9Ö��������1����H����i1�1�����y�z�W��K�τ�]�S�zn�u�w������$����w���y)kk�W#, �~�u��KO�~�j��PV�w�<�������H�X������'(Q�1
K�6�w��z������u{3[�p��j�)e!��d;�ǣ�_���xs���B�أe2)vd �ﴞ3I��K�Glj=�JF�Dg����xJd>gg����/v�O��V�k5�,Eɻ���v��"���v?T���>��o==	#H����8�/�+%��Ï'���-,��S9w�t�?&Π��v��?�]0���`mt��:�Nx�-��2�l��-��Tˮ�"��Z�-�@��g���v+�"�q��EB�k�|���s�u��W�pv�)�(�����7q�3j���EGT���@[����x%'{^�����Dz�")��C0FD��R(���,��h�u��K��(������r�K7�)�5��u���1���+�3U|��9�]�z�i���Z�=���Pq�o;�|&����n2;�Tڳk~�e$���E	�g�z�e��p�����N3m.�C�^����X'�q�q<��V�~t�כ8��)W��멬6,�����
�t����t�ܸo�[`mX��A�T,%c��9���AX�*�wZ����	�mkU�%�̪!����}X=�b�K}\�{�.ɐF���Bȴ���S�]Hךz�G�p1��ED��鼯Y��ʾX�U��چF����q��@��oֈz�ʇ��O�we6��!���V]dJ�
H{�S�H���D�;yٗ�V�X&�݄�+�N��#ho���u�P��G��F7rb���O���29�hA�N��y�6�Tha5%1Q�-#�s�7��}UrRf���1�]�/pLd��U���m���.T��G��q7(�)��æ������mdD^�P�(��!���ϐ��'?o���e�-��e�Q�\��%?����Z̀Ž�n�q���*��1��牆���s�"E=}K'U80�� ʷ�G�FA�����X��)]��x���<EQ���./�:(pz�a�2D]���ݫ��]�?�% c/oG�)��Uj{tP�ތEiL��XAb!q�S������&�c��u�^9�n�<	dh;����]�^ULAm�9�֒O�C�m�hmjj�7o)/��`�:T�����;�d8�$*6�-�q�Ydi�<9����������z�ZV��!�v��zE�ʕ��g�,W@)xrl°�	�|������RP%f �l�`�>�ډ�n�2@^��g��!F�}����A����fTL�����������-�[�Z���\8,dZ��*�\�o�H��2|����ɌTAHS�Ͻ�S��TE���Lx�n	HHE0��dZS�;n!�5��f�4���g	�4ц��dr���WN�(�>���Y�s��Y�>r�'�����GR��On��e���F�}���C�u#��O�4���+�!ܓ�����:�/a�a�D��M�/ͳ���Ed]��H�U��S��wK >W��iX���@��Ư����K��t�fVh�,�닶���L���9κN�+D}��~��.AP�q+'B`#�S&<{ks,��'y!}����m��찃vY����~α���a���*�Vg=������wDR���3.ʃ2���}�h��~�{�:mFY���
�iX~@%c!K���o2i����l�������ڔK`[B�8�h����6)j�G���v@M@|��"�M��,'}�`��Cz�hZ~�+���gz;;PF|>Mћ;"�"!��q1���E�O�pQ��v�~�/�^���D,��pb�Y(C{�{�f�����#����<]��P��}C{7=T�
ʤ��YX������f���C�`�r�nEJ�49 MvU[ͳ��?���J%�d��S���%$�k.�x�,26$��� ��ߓ�U��*z��H8�G̷?�Zl�ҷS��b�)��;��"��C���R��_/Ž���Š�oG�i���=�0
�87�;�x�8���z�9�wW��������4�/ܼ@�T��� ��Y �._�ۦ��o�\�����+����Z]�.���7���PIͷ*D8�at��u�ch�� N;7��.܇�_�UR#\�".�Py�����-���,`��1xCt`�����a����IŨ�y>��R.����K��Zf���P�l����5cd"��`�C�s�;�As�Ox-�b\?Nƴa�|�e�x%ϳ�|�c1H�9��>L*nK]��$A^���r�j=@XWl����q�q�ң�M�|ɫ=:�hy&Y�:t��x��z��\��|1���������kE�VYmE�$X�3�t�
vy�4�%��q�\��`o���yT�Aa|v��p���K����6�2lۜ�ߐ��0�L��(_MdSp7��/�CCڼgݞ���s�Tz�k�e[�"K٠�Ԭ|��EH��7���ܜ��h�tJ&��Z��F5�+�f���1�^ &�9�G����|v3�Up��I9���a��R��u�ޘ���H�S:�g#�n�-}9�t
�Y�4>]�+��d�|l>���=����~qr#�sZ�>c� �>�>�)���U�Zf��:���-^\F�b6wQd�����~�{�n��|5�h�i�h���ĚRzj�I�'��� 5s�]:�z��)R!��x@��)���Y�3c�l������N<@�\-�-N;�PɁXւ��,z�W��� ��� ˎ�x�u���_�I�Rg)� ��p�b�.�g�x�Vyv�G�s�u
3. 	���3
���2�ivtS�UQ�B��%g<�����g⿸�]+��� If�_�<R��+f�a�U��3Ֆ���G�=v�6�}6�!\��T�B6a���xK��K��t-�V_�Ɇ&x%�i���4g��V_4�R{s�����y�;�JK�UQ���!"�[�,N�l�
��Ds�e9�Vq���h0װ�u�ѿ�\�A��(V$�iaU"�.�"]֘�4�Y��y	;J�d���M�_�)׶5�h�͒^�߀,Xw�!\LA�Ҝ��RX��+�`��+=�ȱa���_���=��X�E����Aܚd�ß�<�}��2\T3��n�bN���4�:���~2�n���������9��$���1P�p!mb3�`��s��d}Ǫ?�x��-����av�Z�c�?n��K�gwE��r&�wuMu.�+�%|���|>���0�$��yukl>'`�<dY �#�Yd�����0!�A�H床���#\>�@���'!\��k`��Xjʸ'�%�<g����b7���r��T�����Z�s�b�����5 :�#.��V�Oتg9�#
�}���	�Ӭ���vq�Y�+`\Wc�D P�#'���z��oZ��k�b~�Wё��7�a D�ڼ��O'�o����y�v��0�����-��e���~�X����aZ
G����aL�["<@�b]���(�H+6�ƛ� �	2�lC["�#+����ڭ�m*��-Oc���	��}8F�v;�������V4���Q�^>�M��t$�QU"[�9JC�L��Ƹ$/S�:W,Q��'��&�#c��[�Z�P��Dl��u�����<eT����(;�kY�Q���J��L.� $!>QQU/E��)M<P�#�BKA'���b�������_s�`!
�<어����&wV�]s��"������l��W$�^���R7�Gȕ��+
�O�/[=��ai�e�% I��ƻ�[��]�R���H�8���t�~)�
�CI��(i�C~���T�K� ���vdn�C�B��TO�]�<$>J�/,�J�~MaX��$�����}��\���@H\1J�yN��m�M��~�h�t��p�ۉ��������6�|BSX��پ����!Zm���v�K6����
����rW)�#<�>�p6��lͼx��y�N��/Ժ4�L�wl���>�SePD�p���j��g˯]�C�Lx#NK��]�E*�U�G�ó*?U
:�����sqz�������t�; `x7��.|q\t;!����ށǆ!y։��p�Z��s昏M��Y�̂)���t"i|��no�T�b�#K����n�>XqW~l� p�_M��V�l0N7���S�sM�V�kv�1���j����Nv����	�p��{2�7��k�^�+C��o�w{����$�2��h|!���I����!��j�K.�k5Dҹ��Z�tJ���3���2J�a�����D 5���Qf��L�]��߶�/&�>0e�� ��J��Y�a�����a�Bp͔�ڕ��I��`k�~,��)�>��R���"���WA�KoGBf�T>�?�8��7���7/{�������p�W؎C���ݖ�J	���&42րĔPO���2I����%��&��"|����=��w`���n����<f��B�����+)߿�3��P[��٭ݔT�M�J��q�覱��PA����FӂeP��%�_��>��'��]%�F�{�U-+7�����b��J��5���J>ip����5�Za4���W�-���-Cc��/�{3�2mOѣA�|�&P"�{�ʄ�"������-fN����9�ꨐ��7�<'�����ſ�H�Q�(���%cEZe�_��r��@�ͥ�8��	v/A��M�B��!�����Q�����%?��j��ק����(N�����t�n �|�?�r �X�+Nd<�qM�d�V�l
��+Z2�ݺ���p7j�l�՛�KZ�x��ZӖ�=�z�#��(�T�$B�
WsSaI�a�g[�~j@��P9 {gq\��!��%�0�i����Bo���Q[I��yr�m5�BJ��v�{~��K�Y���|R� F/����7B;g�Vv���s�ݺ���ʝ{�/,���8�hW#7˷:E>��ժq׀~5�*��*=kՅء��OyS?�
��ـ����+�~����B2Dy�	���R҄~� �E&����s� �G��twO��Sq�ئw�shH�O�:]A�1;�N���9�_�G*�6���4�BX��^���S=B�ƗY�T��|���o%����M5����}��"��N�@̌a� _���>?�����%�q��o�@9i��[���ڹ�G��$_�m^e&>j[��\���-N'�x4�r�7;Z���.G�cx�cE;� �o
�d���m�\㕺-��Q'>��c!�/���^�4'Ч����r��p�`��._��Wj�i#9��7@oJ ��� �ܢT�LӰњ�w\)���@8������!Բlފ9�k�lQ"�?C�1�x�����l�?t��@��� ������%ЉٰP{���vW�(��du�'��LgM7
�q�%�&9����j=�(f����0Z�8�^�����!c�T9/�d=Fȫ�1D��o^?���yY��A��Y5���B����ʖ�4�&���
ƿ�s�WHu�?]r9ͨ+O��c(�4�!�($pz�M`�?JKDK����w�7�s���Z��W{������e��8�V!��P��.C�M]�a�]B�ڭ����;�ޮ�[��)�2���FJR���apX.H)����B�_�z��z�3�2wi�v����A$�˲���%�W���o>��+p�O;�7����,���D8B�%�rS��kզ�>������N�0�k�~��2�2�
��2���U�F��m���d�)#�`t�T� ��f|��w�@��:S����k'�Fo���u�ߏ�юc��`S�qޛe��>| �����P�
���Q[�� n�����j�|�š���5o�e��M~���#�
�C*K����L)����k��;
���c/u�[�ς�_M·�t�+K�5�+Q��(E���m��&C��2r ������5F�\:��~w�Τ*����d9��0�Wtҕ½;�YN	b��1��f'�)���/��GЁ��;��#��5|{_��aB�����P�%i��q��@2�O-*�g�'�;	��2D���r���͠�S\�h^S�|�<��R }~7+N-@��~�g��g�d�04��u/~�h�B������@+���@���o��m�Ȩ8�>�O=l.T$sɂ�|�)��շ���<vچ=���&8R��v���G&ߟr�-D�h�t�R�I޸Jr6�}%k��n��&����gM��
"�9���Ȟ\jJI+��0���]�bK��U�(}��4(�{��~h�3�ة��p����s��	���Ue��9�3[����*�9{�7$����~�0i_�^�hu䢶w�O�Fq��L}n�Uخ=��nQ	r����ID��\⸃�$0ň��
 G��-��3�& k+�.��/���}���j�MTw�CFlV0�ݶ�\��W&"8xZ�����3S�$-P����f	H�t������+���;���A��Ӡ�M�j���٬����b�"���HD_V0D�z�3P��������P����-��`}�c�\��<�Ϝؾ~C��>#1�@?/��G�G�H�Z@�ME�E��U?J��΢�����ڮ%�b7yW�C�~��W: �b�9U=�1~[����#�x��@9�W�
3�ڣ�l� }����f`�c#�5n����� ��� �CQuc��9�W(�3�R���zݦ���~Uօ��*Я2�m�y�u;ޕ��PB{��� �bP��T�0w���]�6;%�����)�����P��A���0���Cy�')D�u�冒ҊX�+�f���Bʸ�]���~/6��5ȼ�m|��[�����^��s���O����S�=�J����uI�wQ;!����}�~��V3"�[p�u�}���"���@���G��
�\��sr��ޮ�C��ff��k�i�V���uӫ���a�>,������Vq��l�rE������ʮ�r#j�$De�6�u�ɾU�ϼ�g�Z������e�c�f���( CF *QF��7�܋���	^�Wt@0c�-?v��Z~��.h[W�W��u�	�=9���	��W���A\'4���M@�����"�r��_� ��ԑ��߰���s�~Ѡ"6ύ����(�v��ҥ��8A��sb5վP =T�9"���H�|�8�pR���"	��;��(�c<LO�R.={���&�����0|����|$Bb�-�(S��ez�Ӹ��G&�srR���������F��8�.?|��b�z�C�bT.��3g���O��h��V�ߖ��i�5�a&��E�(�1��8�c�������>f�B"�D�~e�E��&W/DG	A'�G��2�b鄁EZp����o�t��"J����KxAH���+���ݜU�A_|u!��*C�ߦ�?��e�����ז����p�nVlM��AC�������/�:�?�oc�6��=��5U,> -��	F���ND���f�~���[����t�w�Kldr�#��F��ߕ�H���U������N�dD��4��r}�ͭ��B��2,(|׊;�������_�$F;�N϶>d�����J�4�Z�#'�66K�͑)3�	�Ē�q���0��t��V��B��J����Hq4� ̡���rӺޢHA�a��w*�50C�0ܥ��_�]L�K�`���3��~������f�� ��>g�^Mp�#D@�%�[05:�!ϴ*���N��S���I��� ߔ ��4����xo�����'���Ѹ�)��o�&�pa��Q�=���r�����L����z������S���>���1�F�!�A7���_؜�uNI�=؎û�!���m����0"�Әz�	�f�M��j��*(aq���k��ؘ0�Ov[�H.��Y���.ˢP��zhI�<ݜ���@��^xj�z	��5'�7}&�	IɘD%��k���ׁf���H�{�)�(�8� �F.k����O^�����/��G��h�&+�ྐ����.I�gM��&�5v�P�PA�&���L�/۱{�^��<�k���e�[[R2K��@A����un�c����ؠ	[�A���mF�%�*:��^���-���J��{hQ`��ՕH�S�~�p\�"���T�g�wr���3�0�W{1�2/��X�*�'q��Y��������-.<��P9p[,�u��P<9)P�-�(3a@�cc�a��L'L��D�B:�
���;&)NT��E�8<g"ه$!R�'Z���(3}�$4h��_kޚ;�I��c�TO�t�E�I��UI6�ǽI�<C�	$Ӛ��Q�$���}S�y�3T�*�M%l��ԍ.�v|�E���%�e�R8�ξ4��t�W�Fӿ�������U��Qo4���;��״���v�N�G��ϧ�e���hEs�W&w1�!/ё#y�g�Il[��������G���E�|��hv���:v^�3C!R�ʳ�c�/]�!�,�ߚ
�u��Z�c�RA�8(&W�şS�:��0�v�������{$�9�+n�pO�%&A�\�r��+C��7ݸ���lQ�A�0��q�"�&
�%$&\C+oQzcӊ!Sx��^^u�J�#�#d>�L��g���k�Z�O솖p&�(>v���c��dP�w!�� � |�j~��r�l��'�;��*?x�9�:�3i���WN96q䆄j�� �0g��>R���4{�"��=ZW_���>���(� u�2�t9=C�&�H[�Z,�%n�F�� ��k�Ю�����hm�<h������bm>��Y����Ћ��h�	-y���#�p�B�y�Ȕ�/Ys���u^"��lr��� �]\�ɌY���҇�p�Eek�3���GPz��~������?Oa��5{#\;���.��N���;�I�0~|���ov��@�FT��#{u�}��Vs7Ph�1^�u�J�<3@#�s��ӿ`��c�Wsu���b��|TAe%�*�s駋g�PX��Q_�Q�m��1G��.R�I�`�W�	=�k/��`�d/����A#0K���ᇳ�s�D[/������4����y�1�V��p�޶ٺ9�z�Q���#1��[7�~�KnL&c-�|��k#�@�nlr��L!����P�ή�P�tu$���M�BF�,�qv��÷��9ĕx��n�T�8D�c��Qd�G��	,���Q�l�).����Մ�g�rV{J�+������Ծ�\T&�/A[ٳrm�,-w��ğW�o���}��IA-\�Α�Ճ�ܫJ�m=V.��}1LӗM��7��A����〓��d��^��.�D�VO���j���x�^-��w"��+{I��
f(�j 	�&w�� i_K}9q�����-;����>R���ߎ���b�.Ѷ��7���4B�� n�h�`��X�}G�`��ӝ���Sd�N��F��3�Hy���nD8�����{�.S�1]�1�C8�'���]]�ڶ:�`̢��l�VWJ�Y��'�K�C1��5��\���0��e���4R6WKq��@&-��AQ�z^���>�ɔ;d8^�ŉ�Z���{���b�Y\�q$.����3�2�E�m[���)m��XLN�!��s�!�sa�nL�(k�D��:��|ڽN��T/q%=X`���Uٻ�Iwx�� ��@�����O\v��N�o���<k�~ψ�*���G,��Vs�>�,y�ظ�&���t� �4\$&���O&�9��t�#��,����c%�ҭ�q�E��hI��<SW�èP�r���H[�(�h�ۖ.�(	�'@^Z�'f:��ǭ��i� Ü��ш�n�$R��R��pF�I>�H��,K?�F#���#{����L���"��I�j��┩�P���`s��|�u2�P!Q�������!�rHm�}�M��f�~��5���Cy�xi�?�����y�_�b_�{c]�o?W�[�ҹ;QB.������]�U�c:j.�~�Цp�*F|��f	�H+�ݒ%%n���.�ih��֨��&����#%,�H����JeU5Q��8�Me�E�)�x����f}-�s@ϔ�l2_}%uE�voj�i-<q�5���3W&���(S\p�o<"H�w�R�@;8uG�G����H���sJ�OE�	�J#�|A���� ��DrK���	��e������z:W���zr���u#Z�����=/��-��A��m{ ��#�!}�耋4���q�g��ivG���U�*�膦��C�rr���r&��9��Ċi(�%�$�媨�s�9�
gK>��9�x�
9Z��U�����0F��l��{Bv��i��Ф��[y`�*�V= ��zJ��\������7�})������j�z��1����L
���h��K�Y�Ĩ�2~W�A���������[�6�pi��2��}�չIbA��e�vD��?M�P[/���~ᇦ7���G$x�[5X$z�t���A�<��C���(�j呄x ���i�E�������^�R��o�h�S��J�#{��̂�� )j�XErz��m�O���j��$l��͋R�.F�(�Z��UJ��gK#Ӫ�U�*����naN�r�U��Ϊ׎��[*�nP�`q�=_���:�����УVG��"K�o�ĿQ��a$U��k��������CQ��;��P��$��8�9�"X�a/D��$5hK����20����L�- 6��T��lb��7x(1��d'ڇ���|��C��3>1q���%�Ow����k���=H_N(��w�A��!���Lw[�w(c�6��h�*}�V�o"^�@��&�"��]�|'P������=�R&+�ę0��Hw��8���R�R�B2M5P%���'8�m�����.���0M��BI����^.��/�[۷}'��?�l�v$�L�P5z�5}��=�����E5%����3{L���K�;����i���'�x��C�hy�2��y�(�9�>k��ǫP	HY���o8��4�&v���k�Z�h�	���v�%����/r{�B>�y���ɴ��rT��ng�9���B~�A��QMC��<�C����7����@��1�a��j{\i>��~�5����g�j8��
	���I����ڛ��K��5��K���L�;�T;��Q�F<{� ��|������9b1�U-�_n��w��؏^E�ր��iX@��\�k�@�o��F Ne��L���N�6��:��=���wOp=n�ǉH���B� � �e�%��9����N�~n��x��д�"OQ�'>"Z������?���i����y���A��?+M�J�=�:+��g	�>�!*/=�[~�?.9yo��kz��z�N|[����3�)HFk�z{~U��T���#������9T�]6Ev5_ �6Wp|$�q{Rs��f���q�~�o��Y�����W��C�f�$��� }�c!��UO�>iD����f�ޫ��2y��)��i抇�ar�vO�yۅ�<B'���J�͂p��)�i�u���2�#P#[l�������|���ಱ�+��&i�$�!B(�}��"�j�(��������?�4����&�7�1����U�w�A7713l�h+��x-`��ؗ���QV=�SC��rp$vW�g��o�U��%�]Y�+���U��&�^ZK>E 
��I$��3 ��q��	��Q�:��-�K��z3<8��H����ׁɚ?�>��\�K���a�.q��EO�?bd�|w�8�L��x��z�l�P�CXh�=�Ҡ����\����������1x��p����t��RM�\�BD�G�51���}�9L͉x���Y�SѮ��?�X!�&Z���Ӎ؛��Bv�$͈#�\c4/w���'&�X���˵\g�q�]4�
�*8�������u�{�dc���I&hQ��
��G���1t�#�b��@��Qs�s��"��w�4�nm���`0Gu��ג���8�� �<��?��3eΔkd��$35=%���TUi�����Ƣ�d$"��"}�@��PdI�!�(&WG���X�hzsM!��_�B�>��-�2�	V}塜�������ԯ	����������Ĥ���ɑM��K��ruJ���图d�;Q���v���[�%8GkAݚE�lg&���,��C�	p[�ʘR��5��+���ӛe�xe%o?Hֿ��5��p�����.FT,'�Ѡ�?�&U�B5#.�7��-�+ۢ42�e�h�����yN﬋ ��e�+�θ��i�W�j�j�O�}.d�"�dd��[5*�dMBxm��3���*[J�u�+7'[Sp��&u��w������E���R�>ru��z�%�B���{e�^3FH?��!���{w��\���$6�#t?[,��I���EYOs��$��X�˹]�;�'�g'U�� ���ѨX�&��M]�!9z��������`^ak>���#ss�./ga��%Ƥ�b��:�_҃	t!Ɖ�vK{��BR�%W����	��,F����#m�u�`4��V�j�74滇�}��cD�I�?�� ��R�z��0T�Ӥ.�/B��Or�}Z͢�>�N�D;�R[�)�5�?8�� �v:��"���Z���+5��?����+}u`"�Wm�/m�a�}�p���t��$���iot{��!�Q7�W�<]mH�`���+ScǑL���0���(QTF>$�N��_UBYYa0����w�\�R��#f��c�@���5z���ĝ&`�t'S1{E��^E�]�ލ��Q��X�>����t���7/sw9��"е%M+���?	��|["P�U&�����+H���ki(W�0�F�� �"[�;��Sl��&�Ņ���|y�@�sd�*��`�?�3�pH%ov�3����"��%�m�7�3
�l���(�}���(5���I��2R����#!&T�GG�g*���B�����*3�a`�D�[���C��`���I�"nEoQ�w�������!���^�NK����T�]�Hn	̹��?�ۂ6 ����T B��'h_4�y�\;[6D�(����������:���\ݻU�;d�|�{�ʢ}�8��'�+C�4�>2K����3Ѹr�+�����O�%S)=�R�Cg����dj$�u�a�?,"\콁��krh3?e"���!C���M��s���Ӡ�/ud"��A�~â#��	%|E��I����ٖnS5�� ����+ѿԂ�~:n����67�KS[9mA�%9~�	�խ�+�-�F���	�+�:��.�l�	���X|	�^�S��X����c��8�>�7dZ�N�W���iC�����Z[A8�V�`$���{+"U���^�;q/M��{����,ʍqTʰKq�|4&�Z�}�fx`j�?��'@V�%Q�ӏ�1��B�hO�B���{� �����ߏڭj�E�p�T�5���^���0V����워�����e��e6M�Oe~���,�d�5���݆�D���A+:�$�b[U *�6�
��#hA���vC�Z�<؂��F4bк���E9�ɨ#�_�[ת(Ƌ������}��/q�=���SB��@�Һ��[Tĉ*C9�O����3O~�mMh�Yn�Z�$r�j���2s����`�Å)�;��\�~��־�Y��8���qZGJ��m΁v�D��}���섂���V�����Ӥ�L�
�@� ���1C-3��g.[i=������y����+��NkL��AT��!N��W�ً�W�����ku�rKf.Ii"4L����L����;��$�1��������HۚuV� �oL�m��5�o��	�M��%o^�kg�I_
V��O!�^��D�~?���7�Y�υ͠��4z~�X��K�ߋ��8�J�$;��p��%Ɔ��՘88�ٮ�D��ȴ�~��c-,�����r��w��G�#��XT���I|�l�� *]@1�j^��I�`����q������D�hTZ��-̋o�xΗ�wm���ػH�jx�ލ�xϐk�!�sy���Q���p����ȍ�4��H���І!�����%c��W��N���I8�2l�QЖ�!���f�춈���ɖ�ٚJ_3�.�ѱ;R�{�F�F������EfI����A�� ���荒���g�M�I}"�{_9K�a�@ �H��+ح5-g���u�1���-���>��+X�^�ڸ�A�2�^�&�O�S$p/_@W]s��mU%8f,5e~;'�w��1��n��I���62R�����|xavB&�m�7���}+G(�W�[�;sF��2����]Y"\�V E�`�ts3{%
ʩܭ�L]�KN:a���)�
��pO
*�Ɓ�`zU:��`x�ڨ���2���V����P!�tw����QK0�G(4��\�E�BZ�u1����\�CO�F'�^>����{N��팇%sc^���׾i�eXF�5�wV!�ߘ
A#��8��`����Ί�}푿m8>~�������
�̭��VrܟI��:�CK�=���\srT��е����2N]�hL?�9T9E���9_�
��/���W/��Ԑ�|6/��^�U���7�����5�����(�5e�]�7���1Yk���GNx����*Jq��8QIaĜ�+(����_,8��+V���^�U��K�	�x}�^0�z�n1���lS��Rr�骐h0z�\�t)�9�d�YJJ�UY��l�㈵.%�>֌�W7�]�J��>��|��'��8��	�}��<���in�2��+�(W����!�'{����@�cI
F�Z������
vV�!�>���v�7.�b	��qy�	��w���)\sF��q~�<���bƞ�;IT$z��c
_�!���RK.c�J�
��=��]'����L":�!��F^[^1������b@`��Sխ��K;�;�X�-F׏x����lH1�ù��`E���P�֕?��>���u++%d4lql�e2�$9�g� c��j|��:u9Ew6�ͧ����^�<�P �;�/LUo�D�� ?w0<ķ�NG>�S�  �-�A�'ʃ֙G��Ny�\� ĥ�Ck�=�ۙ�:���78#>�n����n���q���%2�����	�.עP��5.t�ݕ��ŏS ��#��pTE����/$D�k�34|]�N)���� K��9<�5��J��\�X)����4�^2`eLѰ >�ekzYb�ɘ�O�uT\�M2,�.��:��Q�2ߎ���2��@��n<�d~����QP��'MqZ`�'���z
�K\M�3�am᣺��R���;����19�S�TO����AY#���v;;�W18d�ay�$��p]�7v?m#x��kT�RdqcDx&���U�4�c�l���J(��Kk�ۆ@F&_���w`ˊTl6>#�{+����OzVy� t�Ќ��.�69+�[����<�M�M���������J��q��D�	��]���1.U����l|������l�NT]�o��YeL�d՛ܪ9���8JT�}t0P$zO���=�ojV<=x�\>��t`��"r:
�{=`����x	����G������t
B�p!�X���bJh>��33U��TA�(�u���W)����X�8Q�r��[�c�@m2���Q�:F�����|nH�[����-�&D+Bat�~���d��l�9��1#蝅B�֥��t`�6V�r%�ډ��x`ZC^S7e:���=F+�^g�G��i��_�N0�C�������~)��nۘ���?Dm�~:K�|�?5�9���1�_(����on�1^~� x�����L���zX�1!=� _�Y,�Bx��:CލT�lT%�Xx2�� �+����|Z��I�;'��B>d��Q�pP��{^؍�-�O�"3��F,Ş��r2��3Wc/���5�T08�����;�9���^�C��܀�i�:�c�bn+�j>��UE��/+@4�f�o�RɮiJX�.Sz�l��S�:/'����B%�c�ss�Qޣ_�S8�ʤ�w�d�v{3?7'܆�#O1���:u�	ۘ�,�Ƭ�H$�H��*;��t���TA��	mG��G���YԎ�����qĜ�=�V�Ը0?f%*��>_�sKD�\
6�� q(�`]@�l��z(��^S���"Vs�����j�Ȯ����D-�j��e�5�=�
�])��6��OS���1��O�i������?��xr�>-3���Y�)l�
�y��ca���S��'�U���>!�]9�#tl��I��c$3�&�"���ҝ��:�q�N�WE�m��(W��O��Q" \S�b�۱�u��dhq�������"�u	 Bv	z`��&r~�us���l�,'��( ^rZ��/��KP���j-`�Ul�����@b���9�]���=	¡R]q �,��d#�����_����-�M���Rh��5NF����kӊv|�yoF�2h_ތv�QtQ�����)S���68���4���6���p�v%�k�uj��v�^��d�K `?O��t�`#$c���"�/�ۧ$�JY���H?�۴y�U@�c#�&�;�f�_n�3��U ��{p��{F��}�I��!�a�-i=l*^��5�}�����V ����T{p.��q��F�w�'��H����G�Au��I������::B*�*���/��L��W�ꭝ�%�)��Q��tū�T�MVY�Vq���/�f�N��ӆ}FH�r-�OɩYh�Ʀd�q�I>�3���b���X��V�ƕ��?�/d���=�+�iJ�Z^0j��ƒ��vh1�y��p�'_�"�n��w���K�F_�Y�>�n8A�%��ũ�m���V0an�^�N����A��jmP��X�@<:ډZ �f	����ɻ^,�\$3Z�jS�DP<�t��aq��!��[��.VJp�#��ٹR��)k���Q��_di�ȱl�6����{�ͺ֐y��_�zW&�2Nrz��9_h���vLSa��&���ﱂ�zhQ(��~վ�:�Y�[��d�����ޞ�]���L�x`(��7���0��5��p���YRit�2�X���S���i\Zm?��X;�Q�h��%��/�g����2P�8����zf�������g�������|H�*wx�`|��ޚN�E��t��q(����s�Y���w��O��	�x���?���:%�1ւG" ή�Zݯ���f�LI�Y�-�8���'maR¶]>>��\f�E�yN`Ľ�@XC��� �����	���H[un
���Kۀ�^����V0Y�f�C���g��F-{S�r���]�9*`]n0l #�]v/�Θ��(���F�Z�*�F7FV@t�Rv2�7���^��-�C)1�ɶ���c��O���ц`�s�^�#9=|�7�5�S�o���T2y�)]��ߤQv���V���$#���_G?{� M�<Iӣc4iW��sa��[�pKYB�f�7�_-F:�t�J:�?������Q%�|�oB"�[�rR`"WV����B<��\X(bz������s�/�b�sh�f�������щ\�!�-!+����_��������h%\��!s�v�����t��Q������ �����~��ܔ7�J`n$i�qK�XK�v��F��m������l�%��7꒴��u>Hc���Y&aL�2�(���b}��v�GH	��j�gV�U�QF3����$�mR2q��
��p)(Ek�-4s�O�W��h"�Q��pyN��ݽ��]����p
���&�)q;d������A�<�J�y���b*���.�q;.�X+������1Ī���h��hW�mA�!v�溔�����6��Č���ě7E�Y�7ٔ㱦m�M����F���5ci�3%_G0����������U���vq�E�]���HV�Z�9J�d1��`0c���� �U$F�ut���'�ݽ�K�[�r,)�W���{�|��Uմ�z:��3H��("��[��Y*A�3�8DN��*����W<+��E�Y�4�j��g��
�j������L�!OQܤA��J|�u������<��� 9�J�F�C9��H�E��f`m��0�#��_�1�"H����(9�w�,����r�u8d���o���`R����[�N�V]A�g)�$����"�Cu�o��Ԫ$����'���ΧpY��t�w�{o��j�;��f��X5�|��:��N�
��4!V�A��q����k#O��w�5��K�\�r�tT�1�O��1R�9_��l��2�M��T��g��3B�WCO��:�C�-�;O�`��:m`�l$M�y��N���=���B��R}?������X�jPn��'#�9�n_B)#4'����L����4� vI���;k����+�˘B_�
,/h���κ�O�#l��up�j�˫o&�ʔg�5D�{H�T�3���58�o�*x?��'ߓdW�F+x_���)#FUE�ܚ&E�oh��+�>�Ib��N��Һ�"��}.9����;	ҹ0�>J�w0Wc�o�Q�OT�%����0�B]�0/��W�t�-�z��ZY���������W0Y򂁿W����s�RvN:S�*���̀��_4fc�/���\��|7�wq^m�&y�̰-���:�y|9nV���}��-E��-���A%�a��6�$�_����%Nt��$��»Dq G�\>z�� �)힩��ӛ!��JTt�E���{"D�$����_᳝��,��������������p���k����q�v�İa+G�;�^qd£�2寇��[0I��&x ���I�X����Ty	�|Z��j�d���H��B���oԇ�N�"���	��Q"҅ő�����,�t�?Y{�w��y+��~��x\���ƥ�s�d!���W�����m:�/̿K�~���r���(�wkS�ͥ��5������S��e�#��
. ֌�;�+Q��r����
 C@�.��^���
Zb>j+�v�Fu �Sl�p��n庨�j���b��Z[5C�s�͇/;Î܄�	B��t�a��HB��m���:a��y4�E�Z��Ն�i�H�u ���QG�ດ��:H�KH�|f`�7�-�B���.*��>X�	j����̿C�~b��V�.��t0��XG �E�c2@��Le��}ÈXپ�,6��$�խ�:����܉N�(����M؂ԧrT���8Ϟ����(�(�����eM�76� =y�A��@��Y?��<�X$��Y�({Q�	ηq�⢦���������%�����e��QL�-x���b����oF�E����5�=�r0v��;�a�!����.�\c�4�mA��}�9��#	�M�1�#�i���2�묍6�E�<͜Zj[�W��m�k~$,L���[<Q�Ә��s�Ib�hd��v�e���`g�Ū3�1lO�@1�