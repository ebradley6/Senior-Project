��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z��4֬��9�A��;Un��Gh[�����<�#�L�-8�o����X0v�c�4��S�`U��� ik�{=�g]�C�+a
>kN}%]q�]���g��k���Y1b	 ���5��G��r>��T�CFT�8g>ڑh�?��H�&RXA��z�b�}'���mR��z�^��"㭄i�Y���	�׍Q�H�q��"SR�D1et�2��7���������)��M���%�dd���q�1��7�I�ޥ�Z�.�m-\ئ�;�#��U��-�G�^�S�+�sJ[o7���O��=���l�B�:�l����PI>N�bP��t��h�SH��c�����D�Bt�R�H5�H*9+�#ã M/eM�w�Φgׄ>�	/_��Λܑ=���J���}ѧ���w'�ōJ���p�b4c��1S�6�Y&a�0m����_�ɑl����ܥ�=�
l?p��j��Ss
�
�E���!������`�rQ%54a��k걱�?)F+hD��̃�v�W�$��F���Y��Y�?�q�޴�ߪ����A���`�����/�`���04� ��7��O��c)ws�(�4����Qg�2��`r�M2��%�`�)�T|>�_W}���m�ݒ�
!:?�D~H����p�/{R��ףw"�G�D��tSז҉F��Edb�7���&�{�lq����ׇ�d^�H<F3���Ӛ��bAR:�7:k���2d��j�	m�����$.k��p��c@�O��`�)vF�J���������j`6�!6�B��;����!Mg �a���O�S8�~F�G��u;g(�lwNZ�$h0�
��c���7��^r=�Q�%n
���� ��
$�s�4y��1����!Y���ּih�Z�0���Q�t�X�u콮�n\~`Z����'t����4����{V`�F�N��x��������(��/�0`�|q�6U�Mpo��.!2�v���V�_<�XA�;����!i�5쵖�-��<'�;uHHāљ+�lY���ڢ��O��[���&T����_2m�-�(�nxK�;�x2�=�ja���^�[h��x7��|\-�[7�5�-�p�6�	��\��Z������yL�y��"+�Oe����?�,���8�!�������.�ޭ!��8b�,���V��]���h�Aֱ��Nr��V�xA�-rX������z�!����|�(��[�}.��j$c�q)��7�&U1Ф1�v�zo�hԶ��STl�Ʊ��R���_U�4Cn�D�( u�Oz�Q_������~�ܵ�ߩ�>�(��8n���7)+D~5-�aG��ɀF�O�|��qB���r�?���L��C�HwaM����W�>����ŊIu��r���3&����D��H���l�1'��-�K�B�sY��]��ذ���gF�9Ū�!�0Na���G��ɒ�xI�-@��/� cJ�H�*��FL��W��E��$��#Z0-]&t(�l��_і��Zg�\��[�_���%�#�]���i6�ߑl�܇Yّ�0^m�����@�S\b閉X�rdI{9.���|�\.'
Z�{q�J�B����7��P&#�C�.�[���
>`*[����L���k�K�=tؕj������׷�KT�Y>����[�d`�f3�z��6�IO�WJ�e�Q��(�����A ��g����"�:��t`K+Rr����恂��RMP�Bܾ}6BTX|7��Ē��<����#�N�����1+�r�$��s�e��gI�@�Ŏ%�Xz�J��#��I|��+�Ġ{u�/�Q{���`�;+�Uok��z�b\b2U���T��+�]&:ML���a
^�,�N
IE%�Y/�n��4�c�2c�qb|� T�!�<,)�GP�	[���l�����8v=iʆ}�!��o�:E>�ƻ9p���F�o�W.iA���V��]D�v���~������9��8g#_����꿌%��a�0��8�Xm�v;��h�/���90N��I($!4#�����^e�钺��9�kH�|���T��&��W�gP�GDݰ��ǈ��Pp��	�B��%̺�=Skx�d��c[L�Yߌ��~ON��dU>�K���t*l�l�d5ʚ�Ƭ[��Z'������P�ٹ���[P|bW2�ii�Kk�ui��2�����P�S��c��Oڑ�
6?�I���)�~,]qN�"���&D����t��;��bF�=���/S�焧ӈ����nO��i��c�	8?�{��g�@J_��`��r{4���{��X�J1FF����x|���.�?`nU����M��_�{C�e+B��:1�"�"$\ko; қ�V�J���0*4T�:����M>�&%�
�t��zuS�>��}	�6�2Sm���[bS�J�;���M%&]�b��gfq�r�|�@�(�����e&3Õv�~�r��{�݊��#UZ�V>�'��&����ⶐRҝs������c�wOv_P	��c�m�j��8;��߾�v��.ua^�~��a'�HЏM���8���}��J���~R�lԛ`�r����?�2�f�5�y4�J2��zx1�%���>>""/ �o�5.ۋ�A]�p�7���Z��ԃ�v\BȰ\�z�|1b�Ȏ�8�9��	�)񼪘�����38�]ש�����4��������'e�
D,?��<Խ�H��� ���{�y� (Q*�URB	3W6��B#������/b��87`"em�{�ed�-�E��g{�=8�*S����y��G=V_ ��T��<^+���!��xk��D��3à>=��i.�`0�l��!��T����К��q�;��zPL�7�\�Q�k�]�E:Q�@�;��~g7��Rj0��;G�Z���(|�%�۲�H��%�?��G��it�V�p�xToo����l�V�Ø�:��#�b�� �|=;�hR�
V��Ƹ�-#�?�nAdv����ݪ1,%B���2�}Hѭ�#nή#+lJ�%�؝�ش���($MIW�B�����v��N�����>�R�Zr�M�O���Ցz����J�e 3�a5Yd��ԯ����&/��>��ۺٷ�,{���'}��(.'(�]��_�S�xz�!Y|^��}��Ϻm팚g���a�� R�q)�'���Յ�V�3,�����ו�Rr*D���q���ؠ�m̯F=��ۂ��J/=vԘ��'�m9v�}�/v�B��-��P!�'պ��@R��(aȥ`}�Ы}i�$Q���[��N-�n���PLZ5lQ>=��p�I��ylm)� ���K�S� Q�.'��%8Ud�|\=A4�m46���w�*daڃ�XE�с��<�c�C��f���l�iH��)˵�)-:2�.�M�e%����k2�4a�_D�ѯ0�y�&���:׾�I�gz%y�S�_�vu�Fx��$�&}�@�c�-�Pir�5Xr�7�V���Z\c0q���ʋsoI��ut��Գ�%P�)��/��t�9!4j,%�)Hh|��6iV��y����-V�-Qfp&�|{��&>�ʝ@��2�p�����7ڳ���ڕ��ߍ,5�t�6g���
�̃b��Y�1&₋���}hw��&=@�*�d�*?>`Ea��_��#�2+��x?yq4;ؠ�{�}����(��ߕk�1�B
� �{-M��8�9�L�v~E�0WtI| q�R�����~�����k]���s،|.p�塟=d������Ḍ�ӊYQ.zFl�2wOq�M��e@�T�n�4�/��ۍ��<{!���[m�j��	Lzqeh3��H�{���%2��)ӳ&���/"v���E͇l�T��� �9�iDF�b��	��Y ��V��L�:��������N�X$a��!�G��������Ab*l���IX@:0�s�Y9Cg������A/ٖ�w����'����64dU��|����C?�<�������h'�B̿��������2��̀�"�PBY�JU��Ԛ8��Lz(�#�Ҳ���Gd�z�h���c�F�/}��%�845�/�f������x����Һ���O^{���ܼ��?a6i�-[��������,A�V�Ŗ��D�+����DjEaHɿ�K;4X{��E�������`��7wv�o��O�����F�k��6>�!���1�3N�Ge�O48����[��X�����Ķ��4��F��M�93dIƘ���Ē5��lF4#�S����S���XPh��+�R}b2�Ӿ:��S*��9���LS	FK�1��m�W,v�� �8K�]���O��1*��X����nl���ސ�Å�iw�c?6R����"+E[��c��~ �U >f󍏿��3�ys'�;3&zi�y�f|y�䕚Ͽ�/���:���Cv�{h2J�hC��tNz��1+c�"����SU��yw��\�]�T�(����Ө|�{Z�=�q)�d�>m�mB�Y�*�\4%FGij�ð�q�?g6��E%�Q��Fhz�o��G(�ڜ����v-u	CJ���6.4��Ö.G�|�He�gA���C����	>ԕ۾��E���Hr�e��`d�Y�#M��>�4,���:\����Wl��ڿ����ކK�?`G��t�>n�p�� ݝ��	p���O����R���y��t�zԅ>*��,ʈP+uF]%s�����1�8�&v���@k��,dBj��P����>v��Z%�����'���f�U�J��{��l�:x�!%��F�E?A��$�{�=W�r��˔�<��Y`�=u�>*���D�>G�\�
�,C�D�E��zU�g�ú����HL�Bo*4L��7���p�A`��k/���h�#�!�x&���T2��w1��\�����>S��*V�|_A�B�ypj���p�[	�;ex�k�!�.ш�J�]'1��(1D�K|�ټ�):Ȉ�$��	6G��o��������.!�2�E�V���J诅i\(��_��?�Ś:"e�邎��I�y$��A'RHeΧ��d�?C4�Z������ˁ|wN��nG���kO}w�k�N�b=!��g>�4�Ѵ5|�ՅCJ ����ksɁ��^I�A�(�r�Ǉ3,�ť��}ksb�:v�nP[LȪKh�ܫ�w^[� ��J�����~��T^r�sD�8U<�B�}�í��>j���q�5�o�ZԈ� ��Z1x�][�� 8���߭�,^����r��$�_���)�D���8�#'T�C�I����Rةʽ�x8"��1��UD�e��D���(��+rk��~��(�LL��8p��!ԭk0(�S��w�K�*�
����H"�E��������&10��M��<����f�M���U[�*�>������*�}��O%�x����G�/���S�p���N�^��̰,�Rg�o_̈"��"ǖ_�w���&ўr����������L��H��ŏ��ὔ���jF�m�N*��W�f�vl�س��CtT����h���:��%T�P����k'R���p�Ⲙ��o�6�'��{C1��U)~]}P�s��}Hp����Ƣy.�a�L[��fq5���A>z�(m-D�9�����|�2�c��Ǟ������s���YOF��1IF��I�J�	fc2Y@���Mh0j�_� D<h�pj��IK�g���Ղ��5��p�Fs'�[r�3xE��Ī�y�bfuo�?@{>����1��fm�u �t���X�d��EiJ����<��ھ�l��y��	��2M��i�D�����ܑ��旟��[�'-�ȋ�C�.
����h:�@�!���z�X>���z`Ko�W	8Q�(4 �7����7�%�A��!������ǖ����"PD��+?5����������	؛ӱ�Bw��u7X�>��G�-G:�U}�I�F���#	Ak_J���>�MP�迲�E(C"W�.T*!�lEZ:��o�e%�R��C4'�yy����C$�Y7]쳃�8�^s���&o��J��+�~��Vݶ}�B��`]�����	CHT���o]M���wA.[��3?��1�ս���	R��f��?�9G�6���٭"H��g_Hg��h>�4�շi,a����1��~|�����	���<�C�v�9��-;D�(�e#ZM�4AC��Eu�ճceI�9�� c,KJq8v~'�ן����V����32ufZ��5��Kz��[��o�\FI������x;��bd���W9�c�+�h�()E��F�@�P�Q��	ҡ�TaA!�z��:��{wܟ�^��ny����푢��t�RZ��Ȕa��v0~鶅F��ha,C�;+�����hFb��O,
\_���Â��}#����Kcgy�健U9F�/U���.��+{BE8��Ť�$�t.ިI K,��J�V{�՜�Ev��2�^�8"=T��t���v��d+�*r]V�)`�$׶nj}y��{ϣq5�DFu۱����>`�}�m��7�U�0a�, ��x߃>A%.i|en��'�0K���<Q~a�o6�P���n�V*u�M������SE2��t�&y%�Gg��3��*��D]$v��Ah2��(���ju?�v�EZ�
6�-��s	�����K�����ƕ9��dTľ��/��.x"�3�2=�a�+I�ţa��Ԟ�7��"K�_NB@���˥�A��E_���$3����q�
�
�z���
Lpnۤ�?�D�ad_%�L�Y�*)	|T -���Bo���U�B�u^6d�gE���5Fב%�cYx�yP3;��4T@�a��U�!NȞI(j0�p@/�hQJ�F���{R-��i4�[Z�Z��Mg>�g2����6�d���xif�8J
�h�	yq9yd�S����UF��#�Z4I
��w�\���Ǘ��[=�Z���6h���R[zǟ��i���x�sL���>���Ċ�_S�w�E���yy͇S�L��3}{%Z����8�m�����g��j.�Ik��"qc�4-`���h� ;�w��ek��I���-�h�@VA���񥯻����j�.I�K}�}V"u�`d� ��$�K���.S�a���xc�\��o+˄�����b��b�
oP���`4�h�Ky_Wa#��$�Z
��>p����A_���r��p�)ڍ��7|�E��n�=#A�/�w[О�ѳ���vov�-y_K�ݲ�5�)��q�{�b1I [�g�\�'����D�%��luخ�x36�ef��_�L�*\aͳ	C�k�����9I�r��������T�S\�!����X��=҇���5z�R�/: ��0k'�DĮ6*T��H(a���Lc�\�l��u:ߎ���D�K���Ȅ�W��VX���I�S# t$j鄇�b:`��|��W�{M����R��Wa�`"cǖ�'2jT�Ee[1`���1&
�����Y��#l�ga�E�����lȯ��]�/�(M��ʜ%�w��Ѱ��C^�5"1`�#%c#�rۼ@�Ts�[�N�x�|5�k�ny֠�����6����#���3Y;�;J�q�3{^&%�n�
�9�L��/����rK�	9�˜64������H�&��U9�F1(wZizzt�(��(� �� �ҙF�s*��6����z���Rw�O���b��O=^F���I�>3�WUW��6�'�g��4n�+7��iv��0Я=��0���@����S��ÛS<�%��%gb_���2OwAk>|v>�\Q���wƷ����:������j6g�b�����`�;��'���ٵ�=�n�N�6/�6m�丁?�+e�>�Y:o�����mk����+���K╴ �m"`��z#�9sAS�p����(������c��m�Yă\c	��g����]4;�F�5I�`�v33Nc�a��VxT��z@سx���d�==(G�?p�.G�sY�m��!R�lTFwF�@�MĪ�E���X!�J T�h��g���C��J T+g�ye#� ��s{�� �C��y��w���ݓ���,����ջ���a%����l��|%�Rv��&W���ݙ��s)5ڡ=�A�/z��j2��
�9��7vIi�+��G.b���,ү��4;�Ģ�U���r��v��iuVW=5C�d0�߻���P#[�A����Mh�8�@�E.*�:�����R��) o]��=.����8��y��,�,���s#�_@��a|Q�������aܭ
�N6xL���S�lA-�C���p/�
�@�$�97��w������Įv��w�Q�MB/�����,��B,q%w�%��{� Y���F���9TI��S"G��-����޴ڽIe���x57@fj�p��K��w��z"B�>�R*^�H���=E�j*�JJ\��!˪���o�n�ѮJ�����Ť�J���	�P�'��ӶYv��L�V�y�(�SJ6K_��/4�|�OP���?SV3=�d�_��P��vv%�1)p���/	<�B��a�״�ߣH����͹1���΀�nZ��]���8m�g{�_�/�A�P��$�z�v�dj���:-���>�����>���2.�/%1�����������N�)Zy�ۨ�X���Ze��P��4u�J0���L�ϣ�k�V�cPM�6���w jA=O�+i4�/R
����32f�T���L�>�B�6~�VGV���>P�5젩�qa�w{S�`l���|�5���O�s&�@x=5y'Q�OU����eA�F��<P�=���o-�&��H�I>9�J�2m��"UJ�\�m7�����
xq�o���d��=Mp��@�~���)=@�T�� l�� ��!���?d�r��M+����e�J��6`������k��]��]��a��j��ܵb���W�&LpX����R⟜꺊t�Mc�j�i�U'QѬ筸ِ�C���iaِw�H��ϖ�Q�u������W��%���#��~�+��Y�m՛u}Δ���ʈ]��WsJ�:i�w��4&�<������)�Q�����~������"�Q덓�;�q�5^ea�d3�{L�X���f�2��.�JI��Yx���=�3ł��������ocx�$KX�Aī�*z��k�������PП��ǂM����t����A�4@�E�q�d�~�e�A���������}���v��S�*to��M�^(��<K!	%'����&�8��.<����dq���l;Q�w\u��uͯ�+�|�*���s;��2	���tX����K�&9����_ym!�m_��eZ�9w�Od
�F���=��/>�Q=(1�Tn��o�<Sr�Y�"���ċq���>��(�by&�
���u#/��:]؇n^�ĭ%	���Y�PEq�����yd���^S���.���¯�����|M�QN���v�6I/U�L�]"L�Zm��3ZBl��C�����j6�s����>(ד�Q�_�o����oq����+����b�3�^8��V%���RC�cᔁ�����.��^�$L5i�a��t�i���n��_�^Mf�����bO��&Ԏ�Ś1D;aͲ>/��f�B����&n��I�T��g�?��~��d�Hdj���Z�$x����Ȯٯ��	��C�����p;zK�����Y�%	O���%��H�I?|-��uKp��lg��.�\d��ϐ��P��.Pւ'Ճ�$ $yٝ�ֵ��&���5���S������pR�qNo8摝����/S�`X�U^��i�,�7� K)�S!I#�|��؀Le��F啦|���(b�	��k����I�;-����u��@{�'��ˑ�j�ݼ�r�t���U����FG	�����f8������r<��&�<�[ b��$
���;�2��KoXv�Tˎ<G(���Jj��m%�`��"xw��Ua36!�ta�J�DYP�J�f���56@��]9m���|>`<b�frc_��,�Ho{�,3��uRu�Õ>��v>�0���X�,p"e�9�fN�W*B�iy�-�)�B*5G2*n�2����8i���I?��e$ܭ�R*R���:S?[��9�t��8x7:�?��Dax�<wp��;����1=�2�V[K��� �� <�&+��?�z��%��1��؃[�5c�z~��R�I[O�.}|�8�(�V2��"� ^*�ʺ�����>,:��|볗�;y"I���̫(�o���bO�hi�Nď�� rR���ȝ�<a;$^���=��޺�_���G��k�ƿ3]j�(��D>�Ү��s�A�������fe�X1�x�ő9��W��/�1�~�b��:P��C����BN�7bkשp���g�����m�ڷT��IAf���/#jS�z���xB�����t��Z�|W�ϝ+<a���[l!��sm��A]�����W�%��fH�}$b�ݶ�/�����Y�Z�NF;R�����_W8��@_ꯅ�;�"Lk����9�59���{ ��]�qlgݻ���11}�P��Ec�Ŝd�hF�3cC�-�w��lWz4���1�I�� 	��n�nqI@�Ugl���D�A���J3~���㋡Ú��Ѧ� �Q@���>�9�K7���S��T�㫤cW��o�Ayt�I$�&��F�ݥn�
+-�̦E�cV�50V`j�{M�B����>�P�P��<'=��S����0b,rD�P�ȥ6_�C�kzUd]T�i�Qxr,q�<�?G�|�������3��p�G�sf�b�&�eki^�����{o&���S�T	�<g!S!	�'*�]B�����^�X��Z%����h����h?w��G�#PL�[�*
=�#����>[�{�Q���j>R��3�^��&!ʽ��Α��}�����M�Ǔ����Z�><�%�"�}L �����
�|�zS��G"R�M��k�n�o��~�{O��A!|����u��\)�BV2q��U�^o�l³G�2շ%�5xQ�̪���sJ5^ka��;9tm��W�5��p�Ù6�St��yBr?�w8�b�.�p��F���s��.Ev ta�	W(��c �n'�?}���St���&mW�P���h&7�g��Bz���������S�� rn&jqK��7��
kL�P�h��_����y����sT��x����,�EY9^)�<_�a�G���O��CS�)�M{�3�]�y���c�B[��(vƚݯ�[�m����?���W���{jX¾�{܈Z���&a��d�D+g7�QL��Au�W1�ds|�,蜼��t��ռE�ʛ��>j��q��+:��QO��"�~�EU�UF�)%�o$�F�M9t�9���K��p�J�"A�A�0?��弍���:�d����?zxhNQ"��.?7UQ����ui������@�[9��*��%q�+Oݷ-վ1m9=���yț�(axC��0��г�.��m t5��*��-E!��x*8M���ǙD$%�`u������	�}\�2 "��A��?�<�9/��u�m����c�҄�#��0����8^DIjI����꒵�ذ����"4H(O|u����D�Eu�� PN�,�2;��?�>��;>l+�znN���Q�S������˧���F˷n����k0�����2��XV�4
hXّ_��,��gX��L$�b����_21���Q6��`r8J'�4|��a>�����w�I���i���8i��
3U3�&9D��ƣ��Y�tC7/?�L����Y���OD�^�XѪ�F�WPI��$
�*{'�,C
��y��h-�Y���L80{�߷mJ6���H[�B�\���+�L�ؠ|�*>������k��?�c��˩i5�7 ��A~�>�x!��\��v�Q��	(����r�Ds�9��]~�s(�k{^� �_`�"p0Ns���r�!�Tͅ�p|�����0�s�2dj�L�l\�$��i8�n��}�efGf���]���=o�Kΐ���Wx=d�>5!Q7Y=ċ��0Le�మ�B�=p���v�.c֊�#��h#w/��畦�'Z$����[GM��
)�}TW�	�o�ڳ���m'z��T���1�9�����=��,�_*FO��9���U+��vN���'��[�AÄ�ݡ����u�?��8|��ປ���/
|bXA��x[K�7A�a�d:WP:넚g��o�`�X���j���*f��fx���/c�N�Um+at����p%����I�9Tp�& �a�r��������2�yG����&��C�I��r�1o��M�*�і�����
IOB�MF�b!���Y��_��Sj�߳ja����?���C8e0 �<y��7�Z�ܸ���:����Nrs�P�1�s$G�qѣ��S�G�Di�%J-�V��o����'�'"��UZ�,M�ٔ[~��fb%��.�][����)�F������N�]��GPZ�]C>VNh]�f�1����O~F<KY|�8D��0�(a�1�!�kܚ�Rb�<0�4dK�.��m��N�­3��f�բg�0�y����S��c|\eε0%pv>��@���O�	Ά�ڕ��:ې�v.�i#9�I���n�6C+ �qf����]/j}8rc���Ϥ��oc&X��Eԛ3���q <��@���w�C�~˰{���)߯��{n����~ǁ��a�x6�ʻ��t^��FU��p�I�]M�]���� �J�6	V#�.V�k�AR�NmvÝ��Q
��2´��z&����i���0�ƖB���Y>c1j<�J,;�O�`���GM������t����O��r�)�n:ޠ��M��R2�X�y�2�=�M������b$�T���mq9�`���':e?�9�9\�[��չԉ����@jDV�2Úz-c��]�X��V0|�H��g���/x5��%�Ը63�6��)�q���J��p>��͘�r[)6cBy5V�=��)EM��co'���:#T>�m�&96�9d�`!
E"Ńcn9TVQ﫾���Aďe��fG�;P�Y�#5)OAp��<�Q�a&��U�1b����I%�E�}4^h���.C6��X���]��D��[K��e�lB�\̀�=ZR<	�m׾�rׁdS�I/栺��~)�{�/=�����������a�sB��1I'C���bÿ�7��'8׀��b���������A,7���܅^��2y��;F��ը�Qn�R��H�K�H�)�S4��"�G�$H��w�>����.���l�⯺|�'�Vp�0���������\�q���L}yH���P���nCݒ\){�}�lW� f��F!�C�8�j$��X�Z���~�!=�/��9 CJ�pEN��� 9)����p���4='�7a�HDL���'�>�c�k��.	�����@��|�7X-gVQ��jb)�ӑV{w$WA��	�D�g�#(t���dgduM�<��=�4o��"&޾4^<�}��ZD��Mb���G�����m��Z{���,8đ2���A�8����k��z�Y�ʕi(����R5�u_�I'��&��:����~��v[9��&+V�QE��,�Q�A<�m�w�Ѭ��1>�Ɲ��u���2m$�cZc�Q�d^g	` 
'�}��W�eS:�����?>���	�=5�	}A9uW,�3����;3YC�k����l�F��%�{���:���̅/�V�-����$���#N��1��l�6[�}!@�����T��gey�n��2�� �{[����2e&�V�Nmg�J�Lj���@�d7S�h���P����YոJ��;yP��N2j�F�(�h�������k�Q������.,l��"�t:#h9��L�A6{�t���*V-�ȋ�:/�� ��ş�zx��fo %�f�l܂���
"��kY��3'�s�6X�޷|X�����O��
�Y�����E��횁{���$]cz|��z,h��"C]zɸ��3Ĳ4�l�?�bQΒC-@݇����}n�[ڠ�B_}P�Es\�PL�$l���(:���S�l��M� �:E}㭩 83Ǭ�G��ո��`5ŪOy�e�Dv���1�D�S�{)��w�����h'��	H6>�͢_�R�u���
k��z�-���@KS$P(��r��u���Τu�q��i�\�ڤ�/��2g�E�.��J�ֹ����1 h���{�˄����sj���5��L�M����<Bp}���eE	�.9����� ?'��4��JL�����T���+u�@�}�l2�OrDW�	MA_�o�)���V&i/V�H���g�a����S��z'����m��`�Q�����a�ٱ�W�&u<W�7��r��6l��/�MN���"%B�[�ܣe��N=�о����"���[�XΊ�1�h#a!Q���<\��nU|+@ 5%Ν���~y'������}��B������/,7=h�8�m��4WOqaHX�?���-w��7����	/���
���@�M �Ê� 	H�Q���:@#���wr�͟��"@��qH��zW���)=!z1�ض���k�E��o����z:fD��"R�Aۅ�Xߝ�>ke|;}a��}2M3�k�@[��j}�bt�����Us~��C'��� �.EU�5(j��/��9��B	tGR����V�hE�fd�:(�o�6�[��H0��I�����������B�*Jw:"+���7�|����W����N�9���@I��X)B�"�	�г�6&欰$<.CXĜK'�[�B7��(tT��@?�MHi]}4����	���լ����1�YHn�h1����1dܡ����c+����u���(�K�e�j��
k�~���Թ0��x�0&pIq�zw��x�(,�m�e.P�e��3}�8 ����+T��-�A�kȀ��hHb-��R�.A�o��s&��WQΐs`�|l��x���:^�]�T�����Ѻ�Dn��y7�q��@�}8 ��N�G�p7�O�u`�E����]�GH���Z��j����~�n�,E�>B&C����agt�pئ �G���T�%C�!ӽ4+�w��e���Ahu�%p�r"���{���-�AB=0mz��F�J)JhoEyZ^��<,�"M��ZqY7��z�%�i�Ϲ^�q��R�{�G�R�����VlY:,�6�iBv1����}Wqk�l��c��,�3��&W��T�2ubpm�+K�$�0[`"��4�߯i���kC"ڮ'�R�^��A��")��s6���nR��P����F��z ��>^a�&����-�M�W��welV�|/��y4-����7�î�������"��G�%F���Y��}���0�x��=P8�3��VD����4N�_����~Թɑ�Ɉb|�-OW�̒S�F���/0�؋��E��a'���J8���c	�(Uϓ5��|z�f��E��5��kI�9y�4�?A�W�K���a 4�'xW��ü��Z��:��f'L�ML0���aayx�Y�Z��9��D�Z/\#����7Tb̏~�aĕ�~��L<����g��g%��0Vł��C���+��3�ܻ�^4
��X������I�� Ҏ����iR����kV��Lȫ��9a��r�U�ɽy)�\\�p�A���]o
:���4v&\a�5��7ʀ�O�,�dR89(1�͔�l_��ߙZ�i�]�h��LG�P(ph��ߊ�i+UG���A�X�<�<7�8��6�)�sw�}2�DƋw%�
��Yx*I�9V���ԅM=z��>2��1d�!�+��[ P��3`^l6������I]���P�f�l��XlQ�v7�j�O��΢�����%��;�r�fd��O�N��n#���	��d�h�@��ԁ����g�;�M�;y�X�ʍ���y�?K��M�6�q
�����#՞��A<����Ec��YW&��ؐY�&
$�-Nq��	+��.X�w���l�~��P����I6p�d��E��OQ�AH���`����n��A��{�3��Ƀ�D�^�חswnXQ�U�yJ��pgBYО����H����>j"45
���zV��2���o�h����J�}���G�0��KI�G��{�)�nx�qf}�C��td�5���w�%�E���b��ߏ"t�Yo?�s���J{b�]L����9��r	��]Z@4j�S%�FeSO{-�oRd��v> ���� ��+)��(_X[m���������������� Gf᫼�E=����+�}oL��&�#H+�����b�T�W�����h G
J����M,5��g�- ̎{7+Y�Ņ4���8��5+X�2tcn�q*+X�"��[���a㷪d��N����ԈYdԦ,�kF��u��j��cbܭ�4���=���x��pRf�;�����8�b�p3��c�f'����)wd
��I_������եT�ϕf�i�K��n]�)��am�!w�9�?�w%9��T�:��Ti���&7�'��s����ߊ�Q��z��@�Zs�:.GIg��n!��Y���t����u|v�8���Q�O�A}�d�lOڹ���s���F�KG�d�-������!��ܕ_�{�6�﷦���-��V�۠�db���`p���d͈p����R�����8N �j7��u;��=����cLM2�[fvp��B��U�;g]|W��c>2�E>9
�R��*��<#Ѭ�ac<Ӧ)el�g�Zg���!B������ߒ���X�h~���q@��Z�&{�b�$���D�&f��ϒYww���lq�f�5&o�w-JQ�8��)�Ʌ1�y��II*�a���A��?�G��G�(Н����t����Ro�N���B���R�qVb��>��<m$���9���7u%�{�=�J��άn�"�����T8��v9P��4�����wI��sU3Y�lz�V5�`Pi�P��@�i]�Xfi��64�����?T�pg���N�U�}3��s�b�!iTua���j�M���p�T�ȷ�:���9�Y��J)H{��>8~��ƌ��������`ٲ��?�h);������4���rNe�s��/�H����6�$D?�Yl�Vn�����|o�ᡘk|�xu�z��ե��1)�r�&o�-$E�_�DFu���$�`�58慵	--L M����cP��k��T;���	�th��-mf��O��:�wd;�<���f]$}kHm��$����F�=>��5W�Ml��a����Y���!ڒ���
9$��n�U[Y���)�WĿ�PG4�$�b]�]���U��o	�_f!�`Ͳ���JL���8&�p&�gm7Q^�7zO�Q�:�P�ʍO%NѠ����\���������)�F�k�
���g�����P��#��H~=6Ǐ��.^Oڞ]�6�qR<ss���@%d�:2U��>�2��6�s��+LXkP$[�Iޢ�<� >�5b��)�?���^6#�hK#��Ќ�b�5����{j^4tƂ���T�t�K���A�4&�'9���'q�l�j�L����`��|��L,�7�͈�R����v�N쭺�]��%�e?�J��I���^�K�E@s���C��X[�fq�'B��?���4LFp�L�]�ِX�>O�K��w�p�hѿJ�XQ�h~o,<=[�Էh%2��2܋~�)b�l��lܼ!, ��`��>U0 ���ALVT�F�2����^)���)&�e�Y�l� ��B��z���D��Υ3�n%�&�5���d����FdL��doݩP���� ���;����cE��Gޗ� <{c$�D��5�rX]�+~�C�#��*���R�u$���K�!���O�Q�C�5�ok��߯�)��%�
&��>��!�w,71���y�,�G�Z������lQPݱ��C0ҙ9۞�$_�=� )Np�Y|�(�Kp�ӫ��W���!&�-�7�U0�grq�#��:���O_��4Fz�Κ�vW�	$Udd�Nc��*(��L�:�I��`��V&xWN
N*�,����(��Fth.��nH�X�O�57b��1�QI�d.��Y�vڴ���"�Ѹ�/���Yi��*..��u�ѣN�XI�0J ,��#9X���1$�x�g����z5�o���ZuO3�c�:������e"�&t����m&�H�]wb���l]�4��FQ��f-Ŋ.ʓX�rN��=��
q�;k�ڲ�	�����Po��)H�<�9���;���1e��5�1�􆙛|4� �m��jAn	�:ڤv9:��AB@��䱟���qܔG���p�gK�.d:Yn�B���$��hLN�o���yb�<cu�Z�������F��
Լ�ӱ����=�5�ud�f��6�t0rj"�A���"	�APU��Z�G�a{Fƚ��۬Y\RLď��b�u�[�o����������^9�]��5Km��_6&��-���92T����C^.M��;��Tw�[`ب�C�xn���\mC!;�5�ܱ� v�����D�ge.lY�\"И�<�!��h�|��rV_&i�<���8I��h�&�E��^$M������9{�.����yƸ��`�(B�(c�1k�yЮ�H	��c���n������ƷR�n"���c$@O[^i'h� f�ó��FH?Η���Gq�?A�iصi�;m�sa��>�ob�6'�Q�u��.Ҝ����f,X%N��-�h �I�]%m�'g˧��Sq&����a�vj:��whvy�9��^$����?��hF��C�_HuO�e�)븽�DߔN�s3:�Uh��'󝯁D��*P����\��7�G���:7M#��?R�:�5k�O�Cѝ�.󛙿s����K���+t���Ey?ia����q���Ie!����V3+{�p�e��i+�_c�!~&�X�g3��es^9�A��Ǡj�ְ�i�3I3���ܠ�5.�B�4�E�2���Aʲb��_t����K"gE'\�	�?��R�� ��DL�Zּ�V>�k\b�NL8������,�a��|�1=�����x�&�Z�����U®�Ƽ����1l���;�u����&�����Kn;��P�\��Bs��=)9$����b���V�m���Z�7��f��k�(G�6���T��M\\��������a0N��|i�����TB�5.�Τ�v���sړ񘖵>�=��� �y[�6� �9��+�H���o�@%�q����KҌ54�Z��]�����ٽ�^�\����2�bn��7Uq�#��z(jݐ'	���G �3�ܡ#���j��������ߡ��p��7V^�0�;%�Fu�(�Q�:�8��WFw�fi15���d�%ϳ�
,97�^��rWܓ���k�l&ߴ�|����9$��
D����k
���F��k�����W���^��z��:H6B+���|�T��]����y�zir��^�~.��E�a�pb����ﵫ�O�L�֠NC�#Xڜiu]��+����q4Cv�E����g����:�6�]�P��@��kJq��Jx������~f��8ʢ,_�[%,2��Eҍ�0�e�����Y&a �,�)F�l���1��浶�2�e�B� �5xM`��>�sg��^?x(��ҫv�K����7�-;�8��wC�z�?�V~�Q�S�s�B�B>=�!��~�`�X-REq�Fy��ے�����x�,�A^�2���ļﳳy|����6Xp��a4�s=�S'I���R���{���x�d�ΐn)��m�T��K��ԁ�� *����+��!�����?N�H��M|�k�i��w��c�DH��f�y�>�B��h8\�3f��C��v���9dVn������*��;��c�Ff��,^�Y�� I+�~��Fe��W�j�m�]!�έ�m*�=��q����?`p����}�i��1�:����KI Pdi0����-n��� � u�蕝I�D��4����Im;O�@d�ײ���("��&c�-D��3����~\�.���Ɂ�P ��(C��悬aA.6��"�]�Nt��i� 6\O^�O�X��?��4m�D)��ލ`ҁ�,�t>�g"í�]�7�ω�"t�L�.���OV~*z=��C�F�x���Nt������>잍�3�S�E�k��l��.v l�H*�Tf�>��q�[ſ�eK[���t����c0�,[�x���׺F��By�mq�ҵ����[�e#%w]v�g3���y�bQ+���y���M[ȓ�"�f�WU��t��qyuw��"l�2�H�ǏM���lìSJ��0�JT�"���ʻ9�?L�"{��J�GP�����=�ʁ@������r�p�j�`�&�&��(�G�KI#�DΤ�7������#�7l+��ljy_��=��ٱ`��ю�s��s�}��[r# �z<����z�w�QC���;j~S�o#o_%6E+�&+7s.|�Ó�|O�o:Ο��K��џ���,4lO��pdb�P"p'd�3n*]/�+�Q���,�$4@T�X��i�(���}\O��o8-n�Ip���k�h�p��>�+j=U��#.���;E��oc���ђ*#��Z�,�4t����oe�[\F�Od6�X�ܱ��Z!��)�u��k���c�9�Qɘ�`�!�&ȳm��������"#:�5����_oya��T_�6�2�ͧ����(��͕��<�:G�"mB�����k�Iw��O��Tht������:[��HI���>�"�U�%3d��8��oO�.[�U>�B��ܣ�P�YC�խ��Ye�ƨ�ǂ}5��O�2��y�VY��ڸ�s���J)l؁����3�nC,�qTf��͜0tWoN�]ir|�Fd1g��[G�>�����J6)�5ָWB�;/���/?�a��� iC�d�}l�T�'��Y���X�Zx��t�Ĺ�)D��k��C�;�$��)z8�*�?j�]�v2��|4P�H�R=h}҈b�%��u��)6���9��>�{�C�zd�zcW
E��U�ȚQ׻�� d^�]g�roH	�p$TE�=�銄�.#o�b����	a+����n���z���+������ɱ�F�b�2��A��Z�c��J�뢗���8����A�t�
� =�TTlf�����2f��(�9�}��(g���ř��0%��<�#0�~JI;ՆM"����.�<�T��[4���,�6���g0"��uk����aۚ��a/����g��l!��I�X�q6�ޑsJOB� )��B���qYh����}�����hVn
Z�z �Z������_�$1:e�.e�UhsX�;fOO�����>�r��J����+49
tiV��٠HwN�_� .�g�_�@$_k��N�;_)p�S�"YB�����`f��-=�`3`�LYK�~�R��l�(T&�3��/?DΪh%��Sv��wϯ<Ĕ�R�^��$�r�Va���PߕX��D���J�1)����������K짺���ҡ誏⏭��Q�n��%�D��y�ͯm�Rm�TD+ʳOζ̍�b}vno�R5�v���L{!�e����Et#U�h�.��K7"Sp��T������Q���[e�2'�z��~UL%T�U`P7��K��l#HU"ڛ�~w��ƝQ>�Xxx}���w\��}eTg��G����98��V䵂٬��I�k��JYX5�k����e	��`���0s�����şlCjb�sטN��;G�Ƙ�Ӑ����"��R�w�����6a4Fs=�w�pB�O�OV"S��ɵj�=��O�%���J~�3\�C��1�%SOT��;{���29��j=w��ѭ��+���/�����Fbs[�/��	}@)�&�8��͏����֊0�iS{=�V�rեa|`�]����0[{�-b	�<�N�f��|����
��y\����G�K�0�C��V���T�'$�Vu�ʤ�ۂP��g[]8I(��2�Kn�9�z=m�N,4z`�\B;Ge�'�D�P@V��w�c�a���oU��!K���è�Ӏ��C���Z����MsFd��!�P�~
�cϜ�E��}磹��+�� �x�p�!P5(�?����^��Sf�q+��\�h�xꐐ����Y�cX!�K��J?ǃY��_8=!g��э2�8=䉇&��,�����8	�c���?'
�#Z��,-a�4侳VK۶�O�$�v�	dF�7���\���� ��]��$ݕ9�1�1��+�֥�����"��L��C�lZ�[:։]{�5���~�7UaеI���	`Yɞ�3 �Q�I�J����V\�#а)+�^�X<
O:,e��]v����`�b�I~f�彵TaEh�~D�a���U9��ޥ�q��E:z�{����v3���yj�1Y9%i�B����͎��Y��u�w"�ڲ?��N�%(J0���"��}F���sy1:��J_�nD�֕#?�qq"R�����2�̢�o��=CL�/��!��)�K�@r������@�3�`z|�q��)5����k[�z�6�<)/>'#�=x���_�zd����7uё��~G4z��!����}T9]��fZ��ѼU�Ϭ�F��~x�	I�r�􇙠
|%mo���,�b:�:���qu}�P�ŕ}T<r�{�s`a#*���re7���?����p�S9�O�SF`/�����P�#J�#�,�;�v�xf�	�9�ׇۊ��̑55���T~����)�e�A�F,�H�Ro�ڃc��\��;�**��).������d��kEsbo����]G)�a�m$�K�:�G*�voz���i��Ql6yY%p:ʬ!��>�R��tkp�q0a�$Q���������/��w�P�6������]�c�',���C�B��ն'��	�Zr�Q���g�1�~��|Fk+/�W���U��Kq܅�Р�D�^�� IC��8,h9�s��n^���Rݴ���}�`���T��POA(�nw����y�9|�U��*)�����4��gD� ���0���9:���!�ԅ����_��������;o^��$��!i�P��=n��،/7*��$!"����0%�K�Y,��;��A��I�8�-!D�bm��<�腺��˂�j _��̉���A�垫g�P�R_x/$� ʾ��n֫�^t���/h�F>i��(�����Ź��!C.�Ҏ�s"�'C��+��@�i{:v������(�PU�����,�&�@Z��Dl:��X���akF���!��"~��5����Ii��́�i+;�V�nN�Go3,nn��QM�'6��ɽx���)X#\�M��o-(Uyy�3�|!� � 4���'=-N��YM�H��O��w��pm�l.թq$�.-�l^�Q:�φy"h2�#���N��Ua����`�U�-Q=qGhs9��ݫ�ʺT�
z�{hx%�!rRc\w�Ɖ|ԇ"���F���l��w���c�7��YX���dm�8��c��!�]b�dEjcJV�@��+X4�ݖy�v�r٣yLYߎ߅������2�"3��O�N!�V�5T�9�J�}��t��9�*�.�	�i����[�a]�G�������m�!n�-�"�!�p�y�B_�%8��"ntq|N!��S;�M@M<ҫYO�bDǷ�.��K*y��uAm(5
)Oa
�����E_�w��rm1��_s��G�u�����BuL�Tc@0��!�Ő���bu_աh���$T ���7N�l��m��'�z���h:�_sZ���܅���>|1�*l�˚��K.G�{=��y��GCC�i_�M��VRa���=��ʫZ��M���bD㛜P����>y�����&�[V��?;��!x���*e[z>}���s��S����rht���?����?w�R�N\_|�2���#��V�>�K=tמ*��F���rc���|�Ź$f��%�+��vBw��D�&`4��"���37��P�zsq�!�s <V�)�g�zG���:f3"���Is1���۪����F��@��󉚘��y� L�2?'{š�BA$�[�m]�ڶ��G�h-�	�a���ҥ�*B�t))���|y�����K�}��>_j�i�V�0Y�[à�+U Z֌���WU�Ф�6��NxY�t .�`4���LѭtW[����݀�D���:��J���3�7{�-�P��:��7dLe�t�D�Ŧ
�������sVY�ƨ$&@��ʸIY�o�,h_;_pB����w�H�0�JR�EdJ1��:��F�:^�SQtNQ�2=�vJM����ݪy|���#���_2l��Φ�Ƽu<X=�Oo�Lkr��!�r�;CO|G%�Y�Tͅ����ʌ�1����^,;0�("��j�+�K���*z߷��Ȅ_V�=y������o�ڼ�-	���/>^��`�@��`$�;�G��A��j6���H�P�LU�2����)�]yA.A$2��0���:��i�k���1J]��F���2�л�!����B���\���O�=
jx��Y��2�M��	L{�.}Hh0k{���c�XB?��ր@j�g�i�I�Z"���2i�BIo]&������JT���W�UB��|{*{7]����^9�����+ß��/�Y�/)c����M,�)�.6�d2��\8�ۼ��{�X�TTj�Nz:};�V��*���֟0�%<��[}�������3��)rpp|`�"�|��W�_��O?�Bx���C|�i)����V1?���j@c�;�&s�M�|�{H-,o��k�`��vʏ5\,�.S�8~���R�(x"X��J�������C��q����0�����E�-��� ��O~�ڤ��~J�T�z��.�>v�֘���2
��伀����*W�%߭;}��;��j��w'z�L]��k��G%~]@DW���=�=�^N'�#A0CF��!�h"ɒQ��kke��^1<�5I����x?eGKi痮z q���]�w,����x�����e3�Î��y�,ݍ�*U�\��@q!��7_*Ô��4`��z��-�YQ��ѵ�b~ac!���KK.�-y�PA�$]fZ,;v�?����ބ��HNL�y�O������#��B#��	H{2���L�R����:�0Q��r��L��l�Mu;����܅'T��SY��r<�;	�[�Y]�L܄�R�\��g"Ag���\����0�X/}h��]�L)!��,�(Cߠ��40yc�m�����ʣ�B`���h��Nq�V�C_��+X��x��hZ�J�48�V��/�Q+���C��=�f��1ö�!�jV�r\���񾴳��-�V���$� �LE�F�?Ah�j�S߱�//`�!�G��^oVT�[�s܀=���u١����罰�E6ՃA2��i���Ą�z?J�;�X�	&������9Q��$�,��4<QM~gk2�/�a���
��o�R27����N�J�U+ ����>���YDBP�cAD���7�el�!���7%��w׋�a�x|���L��7���ۊ�H,��Br4�D$��w淩�=~_E�9���V~fK���ތ���m+��������=�/=c����-^R>���ͅ�29���i=p1ڒ)g��V�^ڹ�؅���[u��LCw�Ϡ��V��đ!z99�4⺝����ֵ
pt;���(��tļ2Zv����rL�?(�N	q��l�:
p��E�pv�X���V>�=�ƴ�g3�9�� 4�9Eo)��(7��7��V7�/���K�kCj>}�mF̴wh�S�*j���U� �R���:�8�F́�P��}_�-a�'�96D(z�'zZ�z0K�����IZ.k��U0��th��Xݗ��5|�t IeLs�7��4�"#_��v�S�6��@�p��c�� 39wD39��M��s^�Z�}����XC4r�kq�f%�E1�+nf�c�߮0]��I3IGMz�S�(.�w��o����0�Y��HH9d.r�B������|�壷�+I �6�(��Q����@��~��=�"� �B7�G���+��*
ox��1�K!�A5�ǡ�Tu#"a�r�?EԖi�8��N��$:e�F�Z�2*܇y�
��� =���I�����y������4z�٬ڽ8�Qz���<��j������w�}.��a�S�� ���85�~D�B���`�nc}�*pb �<��n���X5c��z����i���V; ����KFC{�g�:�}b�`�g����6]�I^�������C��b��4R����ո�'��,�ڍB�J��ƉEwz�F\;���?e<�I�f��[���jL,N(fJ9(�!h�8�i{'����_+b>����$!���,�e���Li�� " k<կ�j9̭�
�ﮤٙ� �����Tv�ت�z��,9jk�����)N�C�צQ��)B_�T��m#M���ϾD+^ǥ{�}���Ó��,���z�V��O:a���h���L9���,l��2�y\����^3�b���gj���#���3>N�� ���\�KܶZ�T�Q!{�Of�ϗ��S�댐�xK�.��b�����U3TQ���7�;�O�$�iO��6��[��풱��z���5�0�ܧL$����%��%��&Xj��W�oJ�� ��ȴ��A����H-�%Mi���l�B�1�M�n�ܕ [�G�k'cl9­^l*�� f�_�	s���²��f��������[*ex��j~۲�����լ9��s�^���y���e�Hbe��MZCM8A��@\�^|���d��d-���6o�٨��x��(N�k�"ǁK��ƷK��5��@6��.fh�F��T�S���EA|�rI�MO�jv��좝���;v	NiYW�Q�}˔��P��%/�)�t�#e�����O����J�-�S"h5��C�<�o��
[)��a�=���ǧ�����9#U�Sz������jUf�}e>WR26�:7'���,�=�Fw��V��D�zR�0����N���z�g�A��$nJ�T|�y�ԟf^-z.H�G**�39�*�����r�Iy����\řgꇷE#_��VA��4��VW�KTh��\͏�K����_�Xk3�)p`���ǿ��c� �ꣂ6�۠���G��.�Kh��'���w�/�U�w�H����Mog������H�#p,T�g��|���Z�X֌�
Bq��E�yj���6�Sl/�ݙ�����\�XFTkT���N؂j�x�we�&	�������4�`�e��L7�ʌ&�ѳ��=$^���)��ɢ���)E��_�W�l��0��)�:`~�)3i��5��!L��T��>fc�b p4D�s㣘\�MV�� BS����Rg�,��[�����BÏ�/Y$Eb.Gd0up4^�&B\�;�+qS��ј�Y�wS��\q��%�|-C*O��pD�W)a,q�J� FT6�Y$��q����R�U&�ޝ��@o_�sɨOO|��6�{��ɣb͵�^+�7��;�:؆���V�d�d�}��/zcv�|�y�_�h�4
�]"���K�7�"�H֥�#���H|��4o�I�@5eL��P��8F�m�&����37~��������ޭ�C��嬨4:)��D2���]���lj�[���ؖ��&he��!�ڋz��g�����������F**��5;�d��m�i�����U���'�1�Td)3�I�JW�Cp��2�|�v�6%�"�+�y4h�d��P��'���J�"�`���A�oFe/�*H=65T��L�5�.�oU�|Y��K9[��稢�2G��N�������&�4��Wh^�t
�xC.Jz��.�P@9�<� ��QuZ��}�f
Fg!�N�%�mXɒ��B����O��k��(�Wݺ�*R+mL� A�Ԭd�&���N��R�}צ��10�\�/��,�� }|,����I�����u`5�G�e�Cn��G�y�E�����͘�1�݉8�c���&��8hJ2�Mbq��QOr�=���3�P�.5w3�����(�܎��Jɢ��3�L�J�G�u��G),��� z��9l]Nd䆷3Y��m`GX5�11bo}�0����6��>?2Z{Z
��\V,�R7��(��ɂӚz�#�e�?_⁡P��7�ڲkhJlp�-�N����*0)�èW/�	S�QdBXO�G]�?wcU,2 E���Atސ�4�@-�ocA,����+��*|�_E:u����S������*"��#�_� Ύ��e��J����z�EV)�N$�7qS�ݓ��/�y�L�:fϸ�7�;~�� E�'F�����W�նҲ��$~X�jݗ�����s-|I����2=7��o�-w�3x���{��:�'��~T�����Pg�a�β�n;��=���'!��Ow�N�ۺN(Y�Ś���\m�$#
L��Ǧ�U1<\��(���>������=4١^��-�ݪ|.	��eІ�i�_'�޷O	����g��������������e,OH��=y!���E����P��P1|�̎������9	)���Ө������^�:5�{�4M�����շq�i�&�E�.|,�s��ߓ���0�I ��
�X�XOQ�>�y�I�弞,���/zsy��؃6�^4�4�.z	p��x�X�����ʮ��[�E�B7s�F#�[Aк߳Bϧ�4L�G�3��%� ��IH7z�lhK�xz��\��n�J�1�.Hc+�>D=e�4pƖ�Mf������9�U)�S����\��Q	C��n���F��&&Ulj0QM��E�� ML��2���w8O���6N�~���c��\^�.�V�({M�Ёj��0���F�Z��]k�̄��+AJ�O���Z�|սb�� �o^z�a��R��y�ՐS��� ����O1%�&}����f����0DJ��n��
����W�t����N����5�i�N`>Oܱ�j�f���<�l�j���<W�5���j1)7 e�9�r�K9�W�p�V��zt�MiZsE d�j5�"�
�z��7�����	?u�<�Ch�'��$2j=�U]21b�B�8�������
J��(�d,��~��8g����4++�Ϫ%k�q��H��~J</��Y����Rʾ�oi�&6�
��4�89t�@�aȦ��O9�0�ʠ��Ԓo���K)�h�B��ZB�S�Ђ�& �<�z���b��=+7ԇ\bA�AoS��}%r�l�ͭ�N�;��Q���Z�Mr|J�˩�d尨򈫊c襊�����`�q�=���WiQĘ �g��ҳ�E��Ed�.Y���)H���qЙ���� 	7�`!I�gK6�dɧz+W�aǔg�Ax�ķ�Q!�ȹ��$?LC�[�nh���7�У������kj~�w8b��F��-,�5�E���ִ���+�S\��e[�H�m��mM'}�@;�%B/�"W�R�G��y�KX����'�wN��kD�e=W�2Ϋ�o�2�L�
���Ŋ�7��5��g�]p�I������Dԥ_59$*�6�����!��,/����R��lL�$_̌c�am�$?D�A�Bw�� �F�rS��*��C$'�s��n��_������k2�<f������!vLv�,�.��W�o 5sk���2�xϵ�'�e8>�G�� F��6K�0������õ��+`D|Ǌ�1�����hD�D��$K�  ~��Ti�p55�P�G�f��w޻��X�&�z`�8������$�cMs��z�Et�]�U�OT��Z�ƀ_�M�GX�4�[��dM4���['��ɚg'Y�Й�c��g�S]c(��0�Єa,�Y�ؑ�<W��.5��Į	����+Ν�����n�B/�̓�+�*����ςJ����]����Ѣ3�hԟy��X	�K.��x#z�a��&𞖲�r�x?�-��bO��Jޗ��� &�����~vS��̡ ���d��a�$j�6�)�ە�2��irm�-�3B���"�2�nRdYp�/HԻ�>1��Z��5C��Z���O����,��1;�3���QR�%�,��s�d���T�EV	�u3����1<t���������'�1j�{�a@)j*J�_����˪���!��W{�ɶӼk�/�pA�DRT��^0^j{W��*GR��c�_@e}���릾���-�4"�Z6�\�;8���r^����I��g��헳%\Ϡ���kb+;"��7���c9��v�>�/�=M9�.��C� �xؚ�yt�JkF.X<�ni����ȝ���8��g{[C�zT�4�~�(/a���ɈT�N����{a��&�1G�Oh�s����=&4��I��!�m&��+q��kj���g�psY9S:h[�́_Y���/p�����5Qu�am�H�g�����e��DlJ2~��WL����E���ol#�9�D�����Њm_%/*Ю�<ώ�V��!���(3������O���)c��Oo��#�1���=\���J>- /V�n��W쉶Tԗ���b{�9�m��i�kfr8W���#A
q�=��U5k|���ϗ���v<u���1$/yΡ�:�ɖ`ɨ�`[��2�-Z��|4���ߠ��^�������R���|Y�|d5$G��W(f��L-�^.�S�l?���f�Tc���r�0�ˍx+i0PZnmx�_�t#�.�5�<�*ᆲ�o��朙*�ԓ(������y��}��Q08����V_C��6"��Yd0`Ѫ&���U���-y=-
���ĩ^��￿�im�Ȍ2�������|0��ނ&̮�ȧf���񪼲V[4�q5df���͢]��ɠ����uudaEu�����.$����ao����]I,4u��P �ؘ4��r9��5�ZH�E�v	�&����ǳ9�QaW���!��O�{'���P�C��P;[��?Y9`����1߹��Yz_��(��!����d�_�m �C����A�/�������w��*��j��)�ģ�,\'�5B�J�F���sA�U�f�*�� �c��t�I�Ml�qO�,�Gf	���o�"H8��f���;"��o,E{5�����!v��@�<��L�����=W�7�����Ɍ��B@���+":fqhu[zpH��|KA�^�#��RŹ��� L���ȃ�#�,wޏdS1��&��tѠHW7�~����vS�ZmV��"��D !�ɴ؁6c���)L4�E�Wƪ��6]l�����R7"�;��0zF�4�)T�����s���D���Q���X�׉Tc�t�ya�A�s5d�Y�~&
̆�n����.�'YI�� Bs�7M��i{�;/� ť<�y#6�7��|=4(AK����4��1�FL�^�7���_�2��S5�un���w�����������Xp�Yp��<r7�a�2\�=;�q�7���C�pXa�v�seJ�g"I��*la?|
����se�ţ�V{݋�.���j6jSP���%�R���2�'J�Y̧�+7�_�^�b��P�#��X��#��V�\x�lyso谾�r�"��k�c���r��@�(,{@?��oZ����a��F�����8�|������a/�k�|c6q�'�F�՟��/�^����@jOI��5�����-���h�����|[{�̦xn!L6ъ�-�*��Lga�r��#��'P����8%�fD��>�����k.����עbϿ<L�������{W��}�l�%=3�������^�
�-����6$��S`�U����������7س�=؇�'�s,��f�kt��"\a��>E�$��Zp�$��2"����������|���6�>���g<�UN�N,��&���49c�<qz ڌ;"���ݪ 
��fv��V%l4��c��)1i��x�W��|\�"X�Rs������YW ���Q'S"���� d��eo{ٌ���*|<���0��}�=]�]�ɔ�<%Č�:1��M��T��$���T<��1�a���џ��EX8���W����F$Y��<�!�ґ�b:ׂ�%ڜ�]I�������/�v�N��k��.|G�������"�a`�ޗ(�j�ϑ�&��oY`-��ě�:�xh�3��[���+K�!ئ��Ŏ4Xn�N cΕ|��Y�-๣����F��� �W�`����ex� 9���ᚕ���x7�T��겤�R�C?���O	�D�&�k�5G��^���Yw@c	W�+�H ��.�BM�4��l,Ώ��d���&��I���"g�zN��<Q;��atm4��M�
[oG��䐊�5#/�s`�"�)�n݀��� ����L�U���lø�@���T~�;hF2�@(����jjʬ�N����WO�m?�	���ß:K^Vr�����S���N�|���ўFD6�x����y�U~��9�"����d�L�8�Ô�Ͼ�},�Ɏ���02�s������8�I�[*2�X��"�_����9zI�
�Kg�9��V����#�f;,�c��lƯ�#۶o���>l�6|�9r/���<V���C=7<Pa�<�����] MsJ5G�g�����h�8��[��B<�r��X�Ng�	&d_�,���7kt,�	I�H��J�$Q�n�Ez�i��l�nRQ4�B���Y��żF��P�t���=�ڳ�ӈ^�!H�~�#w(�d%�i׃�	&��	A�d�4~A��J $�w�g�Ӷ웺6k%G;�� ��N
)���� �`�jA�,^y8�m
����5�`�S ��#���7�4��3��(�w�@}����t~pF� �Ջ�xEPG49�]�)�CXZu��qդ�U��ex�\���k6��x���Dwk�FЈFQ�L�f����j=:������K���V�W��f�V$��`+X)FS��#���Q?�.�mDk�5�r��2O��ʢ��
��&�#4�D8�v*�b~��A3��)��3A^�a�k�.Y'sx���s�|z:�D��}{�t�K�.�M*e�Fxb!P�n������6Ѡ�M����\�⌴I���J�,59��ov6�c����3(�t���0o�����/5U���A���Qm�DQ�-�r'�m�!����^=������f=��	�4[��\$������ކ)Ba��jP$C�q���"�(��5���4/��!�(M��琭�~�rM���ׯ6��;)���u���j�'@?%�e�AFϧ��%@p�t��,��X&M%^�λ��� �lk8�5�1�g�q�4�r�tv���⋯��hٶ;�R���:��aN�+�&}��^�`׫��*�8@Y������å�-7�
O�!��AT[��y����,���G���g�I�a#0jՕo ���&��{#�fUӵ���E%jR��+-K)�4��Ln3��qǜH(һ�Ҿ^�/>���֛B{��u�z,iH��|�̫J�9������%r��`p�rp���	���(���`Ԣ9W@�xy��/��R]]f�l�)3V`78���e�iS��k�)�
�r�'�r��-$H�ǽ��.%?3��}(��@z�3��zu�`�3t�"F0>��B̷��D'� ��v]��J���m�,/zPݵϗ�eO(Uk���#�\�y����'���R7o���F"��
 ����,]3�?�}R���C���ˤ�)=��dƈmZ�����B/���p �6]U������|y,#�Y-� +�=�� :5�L�9���V����D�
�T�g�ޡ�%J�@���.>n��J���C��586���̍��'P�`�1҅����0�̍
�����ё��#���|z�s�\��6K@B��#�e�^�a�=B�˴Ҡ�.��=T2Vw��YQo�Zo	��Dn@v��$��G`�$j�9*S�.5�c�l8�pQ�wx�7œ��*K�nuzz*x�w0{{������nSã~ν�4���I��&F���i�x:�O�;�����7|�?r�e[)n�P���$�L���9ɷ���ݿ��8X+XB���~�ܳMGQ�'9_�Ds��ᑳOL�	�t7��rj6�s>P�p�����b�G݅
��뼢��x�G(hY��v&�״��
/Ò�HoO��z�4H���*� �aN�w�`R�<9��K�|�c��e�_F���ZS)��v��E����|����5�� %]ޟt�?q�|j�S���q�d�_�њ�wb��`�����1�G��Y�C6��:n�!�u�C����_��P̻\:�����&����o���P �zI�8�
�N"�\i*F�d�@KPx���w��˲��"2���L^G�����		/�|�Á���ם��K,����~�6���IK�8������>����'Uq�U3��ܥ����X-���g�fuE�!�
<�A�zD��� ���ɛ�R��S(R���ï ���uD�$V����}�l$�4��yʱ=�r�B�$��R�ذ/��3o=�¢M9��O��->s�,�C5u¶ynȓ@�D���,�#����Z%�`����]�.$��b���yHk5�7�'n���_�.��,e�����|V ��eC�逺S{�_�=1�j3���ס:��zܭsքP=<΄�$�V &y�_n)b RaZ�3�Z|����g=��/-)��>=�o e���p����k�-U4\`^�`��qL˕�K�)O����-�䦪�+>Q�I]� ��^XV�(��ޡ�M���M57*���J�37�5��DL���Fd�bʈ���FL�ΰG�cĈCȭcM_�ؤ��̳i�=����;��"��$&���cW)����(���I�Y�'����%V�u�+���� ����r���V�����:w.�UT�r���@�<��R���Y�~�[����B��l�{\�	e�<l'�Y�9��N=��Eg�"��q*R�r�G1����`|��q
������|�}��b���kk���jJ�5Sl<=k(bê�Iե�cLW��*dJ��{���s�`�zQ
��/
*���ǩ���")�X�����x�,�[�Ҡ�
c�v��}ڧ�U4��g�ʉ�����wI�C�?".�lկ�W������g=I�{���''���{�M	��|��w�9q��]0Q����[Y�]���$��?���	Ȋ1�x"�p�#�Zl|8T�@L<9B����|���m3��	T~݉�>�RM:=p�;f���YE3������M��	����lch��:t4h�{�\�4�jY@`�F %�د	���×'Ý� ;\9�`���YA��i��]���"��j3��]�� ����)=�h��R��̢��;~#q�����M�w�$ �Y������\tl,���o����+n~�X�[�Hؑ�U�D��	m���qĈ���i��������,ѯÃ�� ���B4�O∶�M>�_��������y8/�[�	yI`�W���6?2�$F�Y�^T!�4�2�W�bS�i"6h*����y�'޶������x���J�O;d�� 0Z���5�`��Uf����v��իTJ�������`i}��J���5h���uJ1[�PEt7C��'�6���]��Â+V����W�6/>fE�f�9r���Q<��k�J���U����x� ��ݕ����;�F�V혫��!TOT�X�Ķ�C��\�A�9s[��-�_�WG�8Z� ��^���r�1d�� �*v�������%ڝYv<#�l ����4R��Z���2�V놹.��ʒdMQ��=I��~7�}=��q7�+����׍�av2��qB�[.��]Ҥ���>tO@[��N�����<$��,�5�Yv}96xغ]�RVS�dD�ȿE�cO�~�Sb�$��diI������$�a�f��Uc�t�M���9���![��05tΈȥB6R�t��p�yv��=���]�'�A� n�Jq��j�&_�g����G�;���.*!��J��.��&�T�2�ն�^ɞ���'嚔b�����?lU�#�C��K�Z�ANV��~J�w���?J@([�jefT���hz��M��s����J��xs�Z��~�er��ǝz�����v�d�ދ����m�9ڭ�_�[���q�c�#�%�C����D���[��U}<l5Z�X�y�Bf�{�(�Ɛ)�{ �s�[@�Ͻ�n��,Z�����5��(Fi*fA`�_ҕT2��9��#�J��K�Ы��b(��a�����'����qq,����9j����%����#����/M���SD˼�m����o�����?�*��1��P�'� ����5�B�$�k���j�O4I^y�;�q�+9���<�sI	7Z{�?��g��c5�Z�O�����>�x r��:{�K��v+�`��6��N�pz���¡��.���<����e&n�_�HA���W�GS�9�0�=�u�'s�3'�4Ub�yX�-�.��$����o�"lɕX\�@��.�7��~��t���^	�vך�����WI�����q�G7�_���< 6=@��]�����6Jp��u-�������=|�h�OB���=[��e&�ϝa�D��ͷ}���u�|U��Fl��7~��塞
�,9)-��BwE"�Lc.Q�����c��	|�N����]��ɛ�:���Z������6�D�n��v����5�������8L̈́y0L3���2d�q�]?�>ʣ1}���}	��灑�߫���x]NZ/���<���Ra�"��n�H�� H43�K��j�AZ�5%D��'�����'�n4��T'軿WthH|wO�<��=�V<����m'�����Ԭ��{�O��\֘�A (vܹ��E�����T+�(�!�I`�	?�Kn���ְuC�G,nv޼�r��tH��M5�B�۴J���S�|cL�S(3YL��:�G��~K�Qڱ��h՗�hi�5 �����Wl|��-#�Fadf!�_?>&��'��^���C��:,�T)y�����-���^oy�$e��FVFJ��K�8�(�7ٕ��NHƔFEo��i.�)?�R�U:䉉E�B������'_���,��=�*��yIC��h�zx�a��~ȼ�ao�PsJp��!�B�����]H��abxEc��+��ӛ�����&m}0Ko�o%���J(Ɔ�_A,$�2@o�G+�C&,on	|A斘�}ˈ����"��=�Ȁd��bo�13�Rd�P#�*b�g��>��B��[k��g��]�@B>��x��I�Œ�kPC/� z��ݒG�%L�S����ϖvú9i��.��sk0X���'��B��hc��� =���Օ���.��)�|(pN�w8�)�)�@�߀(}y��Hwu���?�RB;'ߏ�v�.��7D������U��kP����?�&��z�p�O���ujR����cS�E���d�/��:�z�� �E�d��Y=����h�XI�G����Wu#�����X���L��5�ER�9ra�I��df�m��R�?�}�f^���ڦ}��;��X��9�U]{�!޷B ť6��˥>��룟�g��(%��m^��x[��X�2n��b����&Duc"� ��&��P(]�"�;�1������V_��K��x͵s���3z�k8�q#�n���$�l!P�����c���cK�!���H�"����MR7�q�r%�sz����
�VƏ�PZkt�܎��!&I˩+Q<A�[B�0���#3a�!s�8�����W]��QT`�4b,ձ]�[��/�U��^DF�	A7!�(���I���B���?ق�RrM��8ɑ��Z=!@d��o�T5
�/W>a��Й3��,��vpյ�)�)�*��8S�~�" �[~=Y�ƴDͶ�-�m�-qi����){d��K���-"���DD�f�\�a��������u�Q�׈;6��fh�^���М̅I���	�ɀ����R��T%��:�d�P?�~zuk&��"�u��A����K�x䦙�%l�e3��r���dJ�d6�x���d�'Q=���"+P��pI��C��~����~ƌ(�G:alB�ڛZ�(1�h$oSj�Tak?���+#_߆$#������������Z����^ /��'>e��'+f�Ӗ�3%C�}/Œ�4�;vw����@.���3��<��C���Y�k0�&�3��S.��݀�~apk�H�֬�g��)1�<?�Y�X&�r� QY�iqnÎ�Ng�Z�Eo��^b"�W����iV����m�-���`o:;����?a�����6�2"e;� �\E����?"��(���
`�G��_;�Ky��l����wě���-q���<��S���ǀ��L/�%]?j���6Z�W���V�����&�O�S�C���0���x����i���Pr��w	��7}[ �wlpTP�N$8�RӤn^nG�����ޒ�}US�d��\����p��/��
c�q��h�ҁ��>%�,���N�w]�Sr��~b�+ ~D��`�~�`qc/��ef���#Xl��C!Ԝ�s��h��0n��ƫ��B�x�������m�
b�s�Y�128�	,��E��},5�ND���� v��)efGf�u5�F�2!Wޒ)��M���SkR���,c�R"_{�펏 T/"�j���a^l��R����!�ŀ�4 [s�.�f+�u���6�_���T�U�������77�b�d
��$����q�Ȱ�&&�Bx���B��Sǟ�9�Y�j�, cni���{
�gJ� }Zĕ̯�"rو��#�(؎�~�i*G+�=�J����Ko��|�[9�8��>F7NOU�,9p`��K8���D�呀y�!����w6@q��V�F!o��:Kl����bى_���2�ѱs�����VE��J[W�㦺�T�(�
��Ӟ�8�|SY�|�뵅5��A��vC?U�yI��"���
�H(n����L����>�隦��a�KE���s-�Vd��}�iQ�.����5H�Y�6�uF�;ð���o��j�R}2M<ؤ@:��b�X�'�Ո^WR�.To+MU ��W%��p�]Ŵ~��jN�b��t�&1C�L+�,��T����iQ�?P��)����`����g�ǥ���t�v�N|{cߩ^�q�-��բx�4W:���#� [�Ô��N��?C�x�Y(���"��{h=�e3�J�Y��^I�6�Li�Q���4��*H\�u�L��}fϫ�Jx���R���h�2��P<4��K.�'˔�a�|Z��?:�rq�A\f8�x5
���M�7~�(#Х�����?�e�߻�v��!��������+��9O���S�`'G#��#�4����Y�����<p���k#���~"VR�������-]8�V�>��Y�Q�[�ݘ�~�sn����B��w�c���Em�ߙ$��gܻB����l����<��?�����A���	}H�?m�^ޛ���-�
G��'kyl@�R��q#K�e��vF;Eٸ�8�jԔi`���Wy����p�����RMx@.��M�n{Hu��ba�Ԕ�C�'������=�&P��8��3r,7�newi���p����f㴢I�}�-�\���ٔ�h��Y�хI�4%q~οbÕ���=h���^��JSC'G؂�L6;ᶣ���ԫ�����u�A!�R�g��]������E�N�Ym����!��el? �=��^���X[���1k�&��t���;t=7�\�Qz�z���l �t�,�����/x��@���e��?��k謹���ҙ;!��8���2H�d�B�RuDxeTlF �� �G��E�\O-�Mvf�.8�Ә��g��Bw�Nq��-���2a�]-B0�(�]�zb��aC(9>c�N;m��[�Z�i���U?q}ڊ�/����@����\�-���ٱ&k�i��S�a�#�7ܔ�Љ���<bQA;ࠏ�\B�H�a`�r_A�/�MeN�4�Aw���t�f�u�X�j�����j�4O���/'�dU���4q�*�����	Đ��Y��ZOhw��q�Ќ�f�^��U#�[ޠ����}�e���t/և�b���0�T���gR(V�sw���ut#���dXJ�
{Ն��ۣ�A��Q���+B��c������:i��'�#�����A���>��6p��G��+�P&�P�I�sy�����bGm� ���@�Ey'n0��C� �DB�?��h濗���S��[&�WGɩ�<hl�%{��|6�`){ޔ ���A�#��������[�|#����㓦����hr�O��XڻA�Hw�Qa-%�ݕ�㏮��?��T�!�J���Qޭ�4�b�d��Y�7#�:�J�8;ⷷ?d��f�e��ҹ�4�Jm���:��٫dq� �]���|�S+W�D�@Q)���%��(��ahѴ��5������v��sO�Y>���"X���f�74��}��'H-��8��}g:4�������˳�C�]�S���E]ܟy1y�XS���ox�������$�pp���cɺU�`�(U�q8- ��:�M2O �tPЭH.�A�{�)W
-w���yt$�֬�:��]F8Fh�X�6������|͵�f䇐8�����`宭��.4��İ�Ӓn�9Xɠ^|q3Ad|���j���]�i�������6��f�y����� �Jn>�S���E�+Eݪρ7����O���!m��Ш�!�Fix����%'����U�t��r�1���U�6�J�+�).{BT�!cş�&-��@������ަ�W�e*�	��w&�˕^��
'�i��d�m�b��_�qe*3�֐�L���I���d��<op����1���`̛̩��f�Չ5����$�s)i�&q?\�G�zԗ���*V7�6�SM�b��%�j�ɢ<�p;vM�uŔ�EN�X���Mkۗ�'pU��#�'�y�{ZD��J3U���	|�K}Y�y�E�i1.sd1:��B����K*����P�)�C�HT�a!�!��S_�y�î�[r����W=�O�h?�M�!�<:o�Z��Ak#r�v��6�6%�Kܽ���m��H6$�T��W�N�9�?1P�0I�d˖�S��9,��n��߄(+��H�N�}�p����q��-#�lG�t��q����P]ø�mk���j�ɠ��N+p�0���V~�%0�����Y���+�`2���x�c;�h7}�'>�0>Ny��.�+��j�1l׈��˥,��9U
�ef��=_�co�3!��~E�^�蔷9�qS����p%��f*� ��J�]�[zu�4�.�J��r2Lό0��s�^��U*��2�jbfi�Z{��	�lD��AV�n�!8�)��C�ia�]h.��-�����J#!i�F���q�����K�φ^�(T�"��Ud
D �3�4����h���Z��g���{�uy]���za�heM���8�Έ����'Ĕ)���} I�a�J�iM=;J�����N���E��Wb�XJ�;��I�e/ �L:�\�~�+q�����-�٨�HOn�1�l A'�yԈ�hwe�Mɟ���ѝT�=��Me|IRbu�O߫3y���}�b��O�5~����-��9	=� �u���C�������ˎ�c�ہ��DTq�y]jlx��@��y�C��Rr�@.h�5U/�z"͎Q�Fz���'$6��R����h�<�ͥp0�NV4��?�~>�<�@�]�;������V<���9��b��r�
H��7�����/>3�b��}6�B�[�]�6g�v��)����ܿ��V��h�byh=H������`�a����.������G�߃����d��=n���3R'�-�a�����_�]����I|A=Z���?���6hfi_��e��P-ѩM/��(\�a���E�Z�;#̸֕��~�*��i��f����y��f�`+qG:�����-7��p���ٙ='��,�˱R{/� ��S��)�;�}�<!�L��i��R#S4cꡠ�B|q'��x�2��;	#5���MZ*xP�Z�);i�_�,8��买� �h �O�GW�;�z��5@Ƽ����iM?Ix���[��e�p��K
r�"����uք����M�����U��=����_K^�����ݯ����m*ya�N�-9��i�:�A�\�bT���U�ei�T���p?6��1�ֽ�h����}��++����u�~M��uue�p�>e�[�#������=q��h�f�X�� �e)�@�"���IEH�~�����1��z�#���	M:{�����N��vZp�h��v�Q�{���tTM�� g�Ѣ���J>���W� �s�ᜡ�\����2�r�5y���L^��u�/�t�3���K
0���f �b�/YirŮ&4V�(�'͒�c��|}^>��Y�l��J%Ob=��ƀ�Ѧ��m��w�ϕJ=���tH��ől����Y�Rm�Ǳ�Ns�wA���-�D�0`DR�'X��/���vY�� ��-i17������I���1�z��VL��b�|�Go��h���(_��"�v�����yGx^�vy�渊�)����l	J�
��a�i��Y~7`8�)v��%�:~��:1�4��8	ظ��%fdxƺG�];��k�嚓�+)���e��[i ��~���x9�0�ע�Q�ā�=;�lI��k��Y��}����-�g�����Ky�}E��t�e>��C�p�W��vm��r8P;Ie�~�n�w�����O�%]�
s|�p��d��/V���2jC
J9�n@I���Y�;�u$�_���xM�ù��e�o��/����@bj���~�k���EYn��.��yP��%{&�X�^��������h��o�9ߤ����6r9��`��h:+TpZ��_���e�g����x�pNqEn�q�W!.y����*��Z��%�����������E�{4�޶LI-�i�C��ꈡb����=��L~����w���q�;�Ǒ��=��T���GL�ngt)��jm�̏�+������Z����:����r�����'?/�Ԍ��c���
�X�먒mJV��a�M%�pH�ְ��ʴR�{&�F~�S����Ǔ������^���b�~�~}d'�8�E�blX���5�}��P�[g��'�Ȱ#Źq�wna��
��
[�x�B���ݥ�4$�]x�X��p���i��1��E�M�����|�	��2?fF���	��W),���Ǔiu�iT>F�Wo�qjU1cC����n�B�zJ��;R�[YSc��F@�T�%o%�,�* A,Z������?���}��t��^- �L97A@
�m���> p�e���"���AF��MܮH*�#8�g�M4��D��/e>b-;�_ؐZ�x�P�B��i�|>�>�Z���;r	+�Ȭ(#�þ!RK�[�a�R(<�����ܼ�*e���p��"��ԃ�Zna�������Ӛ|��L�V�A��'�GV1!����ߴzg��;�x�����!|�uIkt0�����T��e�(�O�̣��N��!��X�C�g��.U[X��y��lg�<k� 5��X�,�����h������z��c�Q�&�{||E�@����m�g�p�h��i�9�޴C'�)����q��8�d�y�H�F��#t���Fd����g~�`?6mISx6��j�k5R�fQç�U%(�M0RE��5�#����r������^s2O����*�1�7��
-]���e���q�
��|���"7�,�*������/��y�����x�x�qO-���'\dp
��@E�*&r�x	U�%��
Lr�^�Y�*���G}^����o�w;-��؈�r5mc�^Ӭd~��bh��+�&�L�4[J¯�R_��Id����艮�+E�g7�;f�,��kp��[���8�l�}a��lW^X��sv��*؂�h¶'�[Kե���=y/�Ck�7ъ~�
�K�xX�N��p�g�c��'E{Tk�oR7eu{�`����"eO�ř���SEU�6�����n~�>o��� f�{�[v"57*}?H#���SB����b�#�{���#-�lty�;���5J�8�5u �qJ)j��vS��BZ���F��� H�`��=³��6���-�+d�2�L�~wf�v�+Sa;�9[���؏1�Y}�v�!5��b~
��-b�T�l�,�FDQX��u9�X�ǻ$��M)'�g�vGs(��:�������G5 M�	{�
��Է��JW�;��w���Tٹ٠�9�'�'3VԌESa�1�Q^��Rv��}}֗��)��u0�j��\W+��gM���r
%�v~��h
�|���O^&�_9�~�(imBֱ�V��ő��`tD���/�����2�>G���Xc2(I驩�o�[�yl��N��d8�*���gYIa�A���p6S�>�Ã�jU!M]���sT�����X
�Y3rF]EY$��>���,�o����^-Hr����,͞/K�x�&ɱr��u��oo�P̐��h �r���p�G 9�[�s"+98���O���	�|�~]��{m;�p/�7˛�K���7{�6�dX�����3��Wέ��d��� �7���Ctɥ��F�jV������ӑ�Ł�O���
45o�%�q�W3�,�ـ�T�xh���
�:Oc+�b��ѻXŇ�Bˮ�2X9����=Y
oE)1��g�ȴc�K]R�)&ڱ�Y˒ͻ��]��.��/R�73�g��F#�7U����b�ML�i��]6ww���lI�@l�I����I-��m�{��_�3ur��da��[���\���DRB73U������gB��l��W߽���K\����iW��0V8պ9�{d�0���^�9�:����[2�n��ICEβɼ5�l�F�$3� $z��5F���C���?~�����z^�]$�Piq�a����We���*띄�Ib#����� �/�L�zr���T�K��z�|��,��Ϟ�H���g�!8��l�/sbt�ܜ�d!Jg�E�;�ş��>��K�+�V�T�^��0c�BY�9�}v1ց{ȎyE(7=�]C�ܴ��+�[T���2a[, ��F�׊�p�9��ka�^5�AИ�;/�0lSZ^@�-������c���� 2ˁ�tsb���Dk`nt�YD�Յ%-�H��(��4��9�Sλ���`�����W��1:w���ߊc��R'C]�8�.�Ӥ�&���dʅ����&��pc���P7*����+6h�G˪�8/<�,��b+���#�A�u�_/{)��~�ӝox�Y��Bڏ�~A1�UX>��o*MHN��� �l�����DA�]�W+�S[̈́G2.�f�	�}x�F��J�'X��l���/�u�:K<č ���:ȫ䫆 �b'}|�E��,���'=&65^΄Ù�uj�1��6S�y�lNrc�^F�����0P��B����r����x��� n1���&��=��ɱ
��zT����3W��/3��x�kHy9�0��E�9�)[˨�����^�}�l�Wb!�.@�}y �u`a��+^�E�F�G7n�a��&�{��<O�k��7��_�f�N�.��\�����B���qVW�^Hf��,�zø�<C�������
x�����B��hLx�c�;]̌(���¾��)�v�5�G@�p�9���'4�����;-��gr���Rx�m׿ƶ+H�Vb��,�|M���E��ehV�0e��w]����
�g���ٴ�,`��{Bp��h4��W������o��O����0���cz���m����$ldP(��?D���K��o������+��=O�*�[����M劤�=+�
�X���?���+�M�O!��|��A�*J�b���.�Ǥp	�jf]��hI������b��e���?Z%�zU	� �̏��,��i�%Q��U|���qF��!A'�5�,��i�Z��Y<DZ �5 h%����qKR*���B����=������h�t{������W�H��f=��c+\��Ғ<c{�-C���&�I�U"dv	y:���~�Lz9DW��{d���?:8��Ƣ��@)p�ǖ��R��<�A:�.��b  ��ӗɗ�]ͣ*H�n� �6 m}��:�"6��u�,S���.�g�����I��~E���F��A�>�������3������OH|/�l��m&U�i�VC��y��u�h� {gh��=2#����Sb	�[m��3�`F#�OC�!�4�!{[��-��S}�ߦ�0?��=����$
��&���~�8x��1�������f����²�xl��#g�5�?�y�1a�w؇��a��R9|��-�4ރ�#�(a���y��i�w>�8��ԏ���=`�l��ޚ��	�G>�8/DP���d��؈ 'o	F�`���[��P-W�#frH?�f/}�:�����:%��A	4~��_ѡ��ӌ��pO�tC	\��`�	�DO`�F~J��Qݕ ���H��͌�g�������)x�5lt�s�U�h�a�r2y-���C6����18��#���*��
8��u|r,N�0����	�C�敜8y�M莏O*/K긫ـL�v.�k�r� TO��s�	�&���M���:PX!&7���&��݀��s�<F��z�8��&am�������k'����*唈<fh����B�F��\�����Q�O��ja}hx�c�����A�r�9��jk �t��=��V��*�9���bg+��o�d��Mw�a�����π��R a<5�Y�x���[�
��� $R���J��H�Fq�f6q����
�ZD����|��'�z���-L���߀8^"+:�l�֠��T�Ȁͨ@[���5����1dwtq���J�&���.j�x)Z.�2f"ꇉ��d�'��G|�������%��qY��V�o�������`Ǘ��E���rE�����H��Y�m�����ȅ*�]�چ��������rp�Z��qi _�k��V�4%�7~:�Y����/�Z����rƞw3v�a4�EO���'��0�Q�D
������c�D��-q_��]s�wk2�f-Fr@�	�������[/�������	tb���4�W�ϟ����3�����C ��`�:�˟���#��dn��.cW��.�=�*ɻ�����M�m���u����T/'���-�Ԕ{�;>����?�J_�/G���_¨gֹyA&���w�FX�O��xe�O�x�
!����j_,($�+7
��@(Ծ�ɬfU��5�u�P���MV�Sw� ��2�#$xc���9k�2Ύ�U�B+�Y,Q�#&p P�@��p�����G���h����H�aA�6M�џ�&y�y�ܵ*Zx��#���͛o�$��'����뎄��S�
G ��FX�[.�[���x%�^�Q���~y|G������z�o�hs���/��5@�����:���Ni;���=���Brʖ���9�KI�D�N��u���u���n��×q28�.��fǐ��d��P�_q�����T&�ڵ�O�K}�R�9�h��u�u� �1��8����Q礋0p���S�lg�t��F�Y�Dm�?>�/x��Gjg��e���!�Y9l�Kb�s�ۨ�<�D�2v7�b�����{��r�!�ښ��ƙ��	��o��>����s�sv$�̢}�����TL<�Ts��
����\p~�ү�)Ř�+�A
���2��74��<6�j�e�N�i'�]�̳�(/ʍZ��􄙥�B��>�f���(+�l�J���ɍ���HG�'��_���T�m�a�r����532��Y��q|��	Af/zu&�'lw&��Og$�!l�ǖC�\`x-���-�Fy���>o���
�	Н�z�k T�h�N�Z�y7.o��[��WR/
��lw�6�Pb�����ȔR�. �ޫq�m��QH-O��f�{�����S�J��x!�����3h*5�D�>�v�U�m;�ql�r�۞����ȫ���_��u���^�h|�ɺ�Xu ��r�%cH_L�ʞ���{�BJ��L+��Fܕ5� ��C0����n�8�u)X��E��Fn���4��r���E���K����F6�ja��NQ�̨}`��'ra�K��"\��wًPI)�%Y����٩,4���?V;�Ш���	��t+/��k'��e�rf�����vu��lXS�ԗ�j�LC!"�`��Pm���������7�y�ö�%nٙ_�½Z�Of�m9;=�"�K����#I����V��\VѲ�Rl�˻⦷
sy��H�P��.ߴ�-6��|�-��B<��57��n����L��<�붥pljG��cې�C_�w�"�c���(�M�n�$$�2Q�id�7�N�7�n�T��	�����掁�'�9�S�2cy��XB��*�\L>|s�6�������[��
���6I��09M��猿�GV��#��:?ɘ0 B�������2��S��� �q8>c=0S�Z�f�.{�9%|��|�<�wC��Zp*^3i�Z@��c��|ir���B-9^��FT���,F��a��GI�I>�\V�/�~5*�N˲M�R�>?��$�v��n�"�d�s�HcP}!�4�S8����=t�`���)C�v.2�\>B�����j{i�\��,JH��M�3j��I��X��$ÄV�n���i�.��/��Cks���GI'{���ʱy��dG��?B�X�<�02�3]q5�b�@�;QCY�����Ċ]B~�o�X{�ޫ���]�|�"U�d/�{��$em�O[��C�Q�>i���[�L��&t��#ϩt�׳H���L�ɇ}�h�O�$����{E���°�P]1DjGVI)T����6�ƶ���3i̍�	坵�T>�|��g}������#�sA�>�V�馘2eB�ԏ{pl�9��B���m�=V���NO�б"�[�O����d�����(v��6OR�]����ʚ�
J�|�/��h��P�����b�,��p��G���� 'D�+��A���r�Y{{?�>Ý�5l\E��z,V��+��VwV.�s���,��<���˦ȹ
p�b�tw��]�p�7g8Ǧ�s�\��w�}�������d�&�"�{��s�z��ж��򥳅�R~ ���e��4��h�k����ɼ�Q�l�[m���\�r���j���0+�k��d�Í�6M��>�[�4J��J]��k�!d�©`�J#Hu�OY��4%^]��/���G��u�H��F)�{�x)�<��s�򍟂;<: �΄��t�>7���7
t"��7����#��c���h&V0M�w$�"��e��n���:^�o���3�.����v��FoA�|^9Οd����|5�O����&!�t�8yF�vz�"(� �q�ˀ��7K�!H�y9�UN���DE�Su��?jP[��Z��"L�������b�K�$�r�ȴ��}��24���\�"�1șaC�Zz<����w縭VDg^�1���D��)��JD'�!���y>��o�A�֞�{�x�v^4�{�^r���'��.��������H���=m-�������>���7"R������&�/P�}�5����BRu홆��b�
jF+<��%����7T���х(,OE}']�e{�g"[4͓[�qŅ����"Ո[�D������{��Y��D,�A��Z��H�"�TUM�ԇB���+.!���������Bц7���h�z�:�"#��0D�1��Y�b����F��g������㠂���M�ef�����H�3P�y�e�	��!���������2=��;l���EZ���J��q�*$�x���t�֛�������*�>֕�4����)�9�;�.�U���kz�7x("�RU�B��:��"�l8{���u�y�H��H�w��ll.	�S�3��5`���)��ފ���)��� �,*��?V:�E�1p������e���WR�����?ti��@,�W��s�T��?I����>%�P®�R��K�oM��es�RG���;aA�m�!S��L=,�e8^��ǧݽ��D�%���y5�At)�������L� ��4jēƗ-��q���/���AxDE�l����Ĕ��.@E�	#�(��Ju?l�$��ڌ�g+��ӎS��f#�;�?��!p)�kX�����`�Q���^��)@�K\����
r���9bbtH��b�n��|1�W.u'����{�8��f�'+��h��S��G\���l��K��}2Q���j<]�f5y�{/�2��2%L$¢U7�=XN����E3��_$��I����4��O2 ���U,����j�&Pg-[u�A�z�"d���|�P�) ��p2�1������ʸ����=
i��`�;��b%D�8���^´�G����t�{��e3w}z^�G3	`�Q,x�΄n������U�;f�]MY��㭑Rp�`�r�4p�eC7�pI#�JY����/���4�5�$Bq�u���
��Đi�ȉm���d��␾�;��Pm���z�L��`����HN�wǥ4Rt&Y?�h9Wk�3YB���fT�r<>�G_ݫ�A\�@�AC��=ӣ�i:�W_�NP��O��Qv()����7���9SO�9���n�V>���0n�l@������L㒇L�f��~W�g
-�8���	{2��+��8�b��ح#3B���*C�`�l4;6�?~E��2ɺ�h�af��a��j�s��5����m�rZz�bG��Im�H����g���V(�^�e���iO�n׻���ҲQ&=~������^�uO�:xTth����s\s�����C�eƢP�u�It�:�������M����W��߀5���	�u�s��ۭli������.jМҘ�\� �����[b[���~�£���y��;P)��?s���c��X�ȱJ
J�4y.�]Ոl������E"������vx��5wz�A�D�	��r:���x��|,ҹp/�,�!1'��!��������p�8F��܈�#�����5�>(fj��*����b���]=|U��N���&�Qi �G�X>�C���5�\i�>��<��S�o[@g�Z�%��2��	�6��yi�3Q��e�q��e��0rV|��g+��[K�@�c�vQ��j��uˠ�]`�<�*�D�'��@wt��vGɟ�uO�l2��Y՛\����Y��OX:�a ɒ�6��9�#�QIO����>�|Bb�V;��Q�_�k���u�W@�()Vi�3���p����΍+f�M��m���c��Rj�WT��glRǕV�5�)O��pFn@g�R�݈�T�ȇ����z����Eޯ`��s����_S��"h��a����.i�����Q��-,r�QUs�U�OkE��Z�xX�\u��_�񴚕�-E��+ƴ��D�2��S�������˛w���!�S}mh��F��)���`,���h\d >^��:^-��憵�w0h
�YZ��3M�h}�:#�� ��B#Y[]�
�눋	�4(QT�2v���99yDluw�\��S7hJ�ӭ�@M��1�?��R="��>sH�f��i�.e�I@ $���32����ǈ�j���:��1����|-���O9;^�����q��\K����7�A�GNᚠ��N��$G�_@��z]� "Mtd���y�lπW��K�%
�@>'�	�R�&�Ǘ�<�:�����A���ם8b��@~�Q��"?�n���n]�8�g��1Y�=M1����i����{t�<��j���G��:�R��g���PTh�i��zrin�T<B7g�U*B�d��\�'6m� ì�c�,����SE�*/�*}bi����� ��|9�Y��<�����VVs\}����/���UB�ȳ>w��!Y��J�S���\e�6��z,�YJ�P��o��^��5��:u����C<�Fjwf�򠈂w�;����z|[�N�p�X�a�&Z}5�*�w��'�S^��sg}z9!}�����E�/��D�;�pu'�F.,�B5KG����?�����B���8q�7H����ئ&���	�����"ob��4횎�	3²�KC�t&hMz4��Gk��M�V�%��0�+CWY���'���Li���RCNܖ�η�Na ��Ȝ-�4 ��q�̭�^�}�5r�q�"��� �0Z���o!Q�Mx�?���������L��0���@%ǝ,�����x���-Jx:�0Ceٵ��Cx�:*¬��F��bT��t~�P������������ޘ���(���-/il�ã�/��LӒ���ap��S��K�.s���\��UY�i�sZ�Β��b�JT�-����Ẇg�0�i��>�5�d�'��_8�����W�9n�P���핪N}S\7ʺ�kx%m���1�����ѝ��h>� /`�t��VbC���{��l�}u1���+�H~�㯨d���fwF7��R$��z]x�'[��w�N|�����f�r:Qv��y��EΧk�����۫Ժ�Ȋ� �<��z���;���5s�Odm��ܶЫ`a�]һ�]>��.k�
\�։	̹���$��P��Ji�u��!�ŗ^'TO��Kx�}gQ�G�_���s��U�06L:\l���3x5��(�~�7T�Y�r����k�t�4�!S�۳7곚�hR��cH��x�g��w,�������2Lipx�� jʛp�����F}-.�S:�8*��׷��g�7j�JNIZTWu>=ڃT��=�)�.K��,6J�`��e?�㗾���"�*Sl�SXP8�!�O�f[��e�v�����*Qѣb��}�}�iO1�rS8����G䴺�'����}r�7�*> O�6©H�S���zAoށ��k��}���I�NCz<�x�	��Q��" �է���e��2���K����4�J��F�U|!�ُIg|���b�'C�m���y��e�m�q�	l��[!�\�]{OȪU!��@�)"5+�<`�6���v�~"�`������ �\a��e���$9�,X
����qǂ��Y�����Z��߉W퍍���K=���������D{J�[���V�6����T]O�+�V�Z���0�O�0����#t
mJ��ڨ�78�F���TG�c����Z��;��
��
Or��2�oR\.;#��2	/k<�h���,t�_|r��fU.�g�Z�gOL��n��C�7D�CJ�lc
���X���B�ŋ���1��t����R�ŵ�5��Uo���lQt����I��3=�@8�?E���e²��0�A_�]��#6[��D论��Yb "<6F�~�(��&27�-��w5�g��E �"�^�/���g�7�%W�n�K"� �ʙYsƮ��^s����0��l�����~+[>�R��[�oY�6l�hT�N��j��ܚ2�?��f�\��,)�4����ur�'�)?�X��HP%���sCVm�gi^�'v�!=�j2�3k�f������`�eW�w��"�CMv��	m�v�/wE 6�̴�	����,ժ�����ɴ+����)�p4d��+Q�v!>���r�.�;8�KmB"]�k�N9�O
p���9ϙ[���x����R�`?k:N/���r��%?���	���D,�fM�!c�|��uv,�4�l��U���w����@cc�rX�&<��&��q{bL�iS�ֳ\��h]!� ��ss�°���P��YZ�B`�!���g����m�q�:�*����!(?mLhŵ]��UOx__"@�h��Ma��Qn�������n�_�����;`C��^da�8��"���gL3���A�z̅'��x#�?#ݫٔR�2������K=�R3"��|���^@O�k�"�O� �d��a\<$��#WbJj%�(�H�>S�9�"�%��֍�ḇY�J�B2�������ҁ�{�m�g��_�_F�Sm�s�'(S,9��-�b�c+�ȝq�z��e�J}��L4v�]�Á���1zd�s�ᲴN���.&�$T-���(��;1����3�3bcУ7��ƕpNj@�襛�k4��Gd�w��8��f�����p�~�9�ٵ�<a�ԡ�oK�Wڳ
��L��O/!��PW�����AOK`�e�&�VM�6�a���V����lq�`���������y��k���#NCǉ�*����q��e_�i�����\n��?���i���tI}N:����:P���<!���R��Q*vp�&�/y,��&������퀚D;�@��@��`���D�0�?��&k_t� JwSQ&��W�%��J�K�4IB��^렞�>�P�Xi����@t�����ҩ�#n�آ�܀��ھ��Z��߁��&E2@��u"�$�Ri?�ܾ	�㲁k��!,��Bߚ$(�Do��P�����nYk�[54�uf��� �.�WΉv��:�w�?��8�� ��&�pC�l�F��h�,��a���D���"��Խ Z�VH�V�Y�q,pX�MGߋM=�!]4��od�M��{P�M~Љ�s�0��ƨ��up��꺭x�:�ID�S>T�NR�Oqg��Fi��S�X�������@EXAG�Y�IQs�k��s���ee ��7>K�5�\)W�&0� �ݱH������}�M�ߢ��t1*W��g�!��P��do��j��M�1��_�#�QS�]������0�Y�
IY�[�8�Ogp�sڳ���-&�a�}�<S��Qȹ�}��b�1n�**zrE4���忰\�e5ڡ�-lV�7��\��J��/! �|ç����T��'���������+�Q:��F��ea���9�tR6����J�����i)�~�}8�����Z�:�l��EM�Ś�����B��.(P�C� tU�T�E�\��]Qɐ��?�wF�8�f��
�;��5���0��[��(�H�k��������ОC^D��K�������C>�л�������>\��0SY��$(��+:��d��Ii9�>.T��l?M۾S�#3kK�3�����_`px3:Z;3m��v�;�(�UT42�M�׉�G�_/���^��4�c�6��HJ��(^0�t홫~|��;��ʽvO�dLL_{K�¨�-"R���~b��n~��(��6[➽�4��ڣ_��&�[M��byu{�@n�g
��!I��A#vᷴ�whp�_�One�τ�����a�[�|�}�̛�	_g/$Z>��Uh�����p�Tr����Cҵ�sF������i4���}Y5-��xiF�L.�f0P�\��d�Ж�_���l����m%�Q.�x��zO��;:�Qr�6��Ire�"h.�W���p}�����X��mF��p�u�c$�bb�8I.�'���88��y;&���>G�:ڋ��b��B�! �sa�h�;�Ƞ�cg���3Ě���Diw7�W��Iw�ƅSFݛޱ�g�t��B�e��tQ���i����-��))?Ӹ��[@2��dqVU`�3v�p��pnޟo~���5fz��ŧg�$��F?��L��6w8��!�IF��9�Άp�j w=q�^��'�Z\��@
�|�>��ۏ��*�_�o�y�2�~���/�g����s��~a���z�(�wX�pB���7װt��$b��liw�B��0�gQ�EwB��ᴿ$�g�GXr$����.�0�n��[�}D\��Ҹ��kŅ�wz��p3:�-/��TDL�����@|��w9 :f����H�~{+�l�f $�������}�(G�r���S̯�%�Ȟ(���R�Y�w��D3����/�?�(�׀��+��$h���Rqqc��Kq�׽�7 J����[�kᗦ�A��B1ѫ�&x�
��a�|À;��ITQ�A���r/,�q� C�е��sk{�������Vm��mb�O�f	���e>36r4eims��=����1�bț�w��k�P��a=;��cH?���ɘ*��O8��q��7��������u�}E �h�Rnb��^n��G�eʜ�c+(��`z���Y���U�AU�=kN�<� �+��'��]^4��Y�����0���-�R�M�&_����� ^ ��`ϟ�`n�������$���}�c������X�M
ٳ�*rԸ�/���J���:Ǝ�Bú�>���w����ɼ(�oAN����|��t�H���-\{`(��3����pp�.���ߞ���<�j����1�*ĳ���fʲ�.P��Vןjo�!�B�)x"_�bn	�x��I��{���$��j쐾�����E�<�9!5���3�����}+y�%"0�'�����S�j��؇��lS�];O��������z��r6|jKl�i�|�+a� �Z�/�*qF�x�S$r�f_�]T�ҥ���gZªj��3�(�խ�����SD�� �}s��*SWV0>A�S�w���a������a[��Dc�WJ:���f���Gù�ȃ/�`���B�Wx�@�0�cfb{�5Jy�X
������݅�慓�vqg9d�r�~�9fvM�e��f���`\Hʘ܈�B~��k��D��;�5IgO7,�uebӨ��T�A_A�rF�Q)Gג_`��V���+diM(��)i�]MȄ9\���*D��+@E�]kiv ��?������a�c"��Z�5�ɶ��CLxR�	ߕ�3�l.�O�.�u�W�&4�i-w����]�Be�a���)�Wxo�3���[�x�%0di� ˗-: �0Bn;��W"l�5(Z�|�2�R"^�6j�p�&��8t5��w+�D��׫^�N���a`�[�^����hǱ�|:�UiNP��nB]��NwU+T.+��֩���yd|���-� hԏ����E/� G5��^�ml���O��h���W��)�� &3���}�9{Ъ��������h���*+��J��$Z�^�2@$
�%�6��IY�<��`�cyg�)L$�oew���g�z"|�O�Ž����(�z&�V�]+Hֳkv�O?������q����A`k�`^�ۘ~��#Ò�~9��`*NE����X:�'��S0�[v��p��$_.U��/W�Pi�E�?��ӪCM�,M�q�zȠ/���r<��Kct��ӚI�(�|���M��;�P����r�/m�w2 �'IB�ͤ�ȍ�@X<+�|��e�lb��oK> ���ϻu���:꩒�Ā:BH�"c!Tj !���3���F���1��/M��(	����������o~�4M��q9u�����	d�Vp�ǜ�p�V�˲J\�-]�$��#��e/{	fO�����j-�-�+ b��~dO��'JF��Uz"�; [��-��t�����,��h�;�nBy���LAɃZ��C>ކ����OEv��p���NQ����?�B�_�[�7�e�0�̵^�"��:r�7�Ogux;� k^9�#vq�+��cqm��`U~B@ �3Ҙ]�	㤕��]C|>y��DS�".6`�Ό7}�Wl�h�����Po��1���o�X��� ���A�3Z>L��W���[>��V�1���\S͌��
5�4@B^�{ż����[7��|��̢H6���.�ׁĲ����CE�-r�\D쩛+J�+��p�ԝ�G���"�Gk�t*�/�J$��@P�������_�/�b�Жo���T1�+BNet�)����;]㏆ ��Z��H}��\4�1Ġr�N�����1B����
z~���P=Q\��79�ʚ�cs]�ï�㾽����z��
uz�������.��������w�o�u�{!���
�a��,�����&��2?.>[�4��	GA�TA�HMA�Ѱ��`W�[�§�����}�#4S�V3{��P9��`�dx�t;����b#b��ч�M�E�ݥD�?�+��x�9
�9ǹ��MA�9�<�1!��T� �\����k�� eL��C6-��7���f�|���_u���h�8�%�_�9:氋I�v������;uhv"����+zl�Qc�b9�����$��[�T�K��|kW��Ú���B�2�ǰB*�!l�3:WFe^jɪ�Ztʦ�F�	��mI,S����Ru��8
"&�	��y�q�����{XZݠ�+0�D��0���`h��1�ǂ�NO�cL)�ج�ơ�E�k7=�T�Q����3Ú���k%��0�*˚���	�	��
�[�kj,9tܐ��F��}���e�u+ ��YEP��#�Qǫ]��l'�5��aܷ�p������D`��n���y��|���d"
5e�f�����Dli K>�:�_��\�כ3
m���W��fo���S�{�\] .�d�x���3,BP�%�QA����ўJ���ْ�x�Д���vF
�6ڔ�M�^Yg
�*_䣨Mf�Q	H��V,l{���Fy`
�a Q`5��=e&s�#�rZ�4O�<���_����|j t��>(�����h��A{�gk<��I
�Ín�AuLi���.��4�˰_A'��b����G93Ѱ��՗/�:'(�B)��Ki�Q� ��\��O�<?l�g9� "d�M_�f�_��$���l�le#����lne���J �̇�"���z)��|9�i�kRw%�I}����0�,i��L����Y3����:,+;�*��Q�s�wH	{z��q)�0��Ҹ���!,FB�ۋf��.۰i~�������A��x[H�'���0j�j{�2����w�4�Y��:���W���y�}���(g�����J�L�Zl�/��hs��#&5닰G����xk�}���0]�DZ�% ����ɣ�D	sWD�}����h�����󜰋y�h{���}ׄc�	�.�Ǻ=��5h ����P�թj|�����^��4�| ?岎>�K7/RS�x�(�LR�}kB�RCm1�Z�	�&�{t$��u'S�v�������е|�ə����4�6�n���ۭ��6�	�5�����E)^)��EXYK�Éd������Œ鿔�V;�.ȧt$R�xH���Wly��;6�ނ������1�a<��0)��K��d�D�#���V��W|���\�XWj��x���r ��x==%e��^+|[�rr9@&�R����R�w�:�^<����N�?YU9�'ސ��'k(K�Aj!��-��*�.��&�����z��F���r���*y0i�����/��3C�Q*Y-$�9VnӍ� ��yڽ!s4��	S�!p�u��3�d�7k���N����V�H"0/$�>�>�����,
tA/F����01�?_w���0�(-n�CP�Q��|1��I��Z\e�D��y�v��2�ꖍQq�:�~C8֏��JX,?BWG>��+3D�X���?�0�~~V�9�����"�铭�t��B{J2n\�E,{#��]�r�p�d"9�*J@xO)u�Tl��H����n�����ⳮ��	n��#��3��[���P\�+O� /\���֬P��_��I{�X������J��)f�9��u��D�yv�A�5ܜ��FǬ�a�7�?��^�d�s���t��]_�1^W�H�Hi�N��B����b��]��}������y-�.I=h7�ld�˛��d��E�4jSE�<k{�k|G}�tMf�����6?�q�"sw���F��ͤ۴�x���%(��Qu:���w�ͦ	�:�s}rO%��K,5O��?*��'J)&���P��r.����9��5�@Ԏ>_F�%ŵ�`��]J�b1E���6G��֐^�K�"��z����M�Qw� �E��9�L��8ϻ\�����,9H�8�	��c�r@��Xb��BL������()w�)���-M���q	���U	_�ق���#��BY�,J��箃=F��i�R�j�B��5H�$*��D���NYկ\s���|�EWY��+�2^��Z��e�M
��&H�ɿi�wnЃ����m�TV�[�*~�L��+-��T�lGR�J��БsA^����m�2WX��,�����Ʌ ��yyv�M�X<m�MX�\C��:IG2�WFl�5X�-2"���������6 �+^&V�!e&��?���M�ɻ-������ɮ��X�:���.S�� 7%���E�.�����U��ԅ��Z�c%�!S�}��(�)�<�̚��E�E��9,Q��&+������9č
c������ S�||�����1������	U�m��V����p'r,�� b���;�ݵ��
�	5u?J���F���Q<�0V�ӱ(�m<#>r���W~8$K�u�ˀ�+E��a���2��Yi8.>������OW�{:)�T|S/[�4B�֧�i���F��|
q���yG��m�;��H+~�z[�D7Z>;���C��t>d�ϑ��kQ)���M5�)ehS}2G�]�P��
����^��hNr��q�ĉ=���+ �w��.0I��d�i#�T��e��AzK��O|�������G&��y+�2?�4�H��k4{h/H�5k���	_���H���L��JI�Jd�Hת��Hq-��0��B~�C���K���&���������|�C���at��ZP;��٨���!�G�62-�<�%��M;���5�l`3���n�A� WՓ�)h�� !�δs��b8�Ԕ�ė�I�j��ML��?!��әG�/�R��
u(�����3C�c�ۿ�镁�]f7���]�H�V���K��e2�M����H~~��[k�g`*��+6�[-mnl�A�^�H-	ل!��� �):�k�<;����n���[������S�_T�)��h<8�l�_n��}OL����4$kƻ�Y�ɾa��"��������roMR�zP��j��q#�2����*���dH!�,�+a+�8j1gf�k�>�$�S_�` �ߝ�e�VSU��b��A��r����?x��������U�?׆�,"ߎuI�<Ґ��і(M��tP����EQ#���J��
]��7�Kt�2����}#�)%�����xX�O�=⨨ w4efD�|ZF of��_Cu���"�'C�P�s��GRWD3�@K�����OB�V+�8>1=��B��D
^�(}�1L�f<��y(}�D�#*0�z��6{Q%�O�-����0�(�@������[W O)��A�q���j*��|(��r�U����)��� �[ŗWAsf���������Bට���'��֬K��pq@�1l�򣋺ȫ�;�w�7��R�8���I����"���b_s�s˛ƽ˙�G�n�ϤYH-�4��W�o'�kې���QL�v�W˅�X,�^�������'�7��	�/?0ћ/ް��{����_Y�vD*I��$,p\`R"��E��}1�v�d�A�S(u~>�$��W���Af(y�ō�)oN�����F����.��à�����;!ֿnI���tE� �?�e�팒e�^�'㨭]+o��Z��+���� �
f�}����z��Գ/ d�ົ���x���r)[I��`iu���~�2"E���̷noP|��r�v�eC�'�<,}�������)�R�.g}��=��ʴ��3����h�[�a��0H�K�\P��c|�j�<�C#3���-��nqwC�l�Y��Awb��C�߿��B�!PDS׼��hr�a+S�.҈�s������h�U͘�=dnm�g"�.��%i\g�H�|"�Q��kHy�1G���@�]~�o7�_��3�"�Xs�|�5��S��sӧ꡻D��'YI�&�>|�[��:�z��q��ӊ%r�쩋49��w_�.�wX4���?�E��!��(�>�N`�L�r��y00���)��4[���W�@��)��!l��Ik �/�r�!�۪����bc���~�����6���O�8��ooǵ�G��F�:Y�<6�"Or���ܒnO�F��]�Ki��Df?r��%X?�� �K���^�`����Xh�5�7�@���jo�,�8��D9`~�i���%v��*�3f��e)C�:H���J���Pr�
�J���\kgb(���1�O8��!a6qe�2Ġ��c�<��
&��,N;�另����4͓����<��3������OtU�`:r�/�- �:羳�D�<���U[�D�W�gb���b�8��oic�/"�?���uA�Z�jN3�Wg�b��xs�K��qX��U�W�Əa�0�����m����i�{c�2�"d=p���g�6�^�q���TS2<B��k�}�G��m�9�E��ܻn)���B8�/*c��O5q��#�mu�u�Y���?���c)4g.�����r�'>/�7
Ti�~�����d�ל�!Z:�&Ʋ��RL��Y("�C�X��+ct��1�f�z���ID�/)�I9���g�`Z�<B��S�.J�O�j�8�bΡ����Vd��*Uz�+aU-;��Ԉ Cs�p�k��d����D�"A��Ϟ�I_ :��J=��P�Rzr+��̬����x`�͡O~�L�b|�`��9���&Z^�Y�э�D�Ҋ���T�,)^��I�y%�:�U%m�Ł7�*N��`Dl4�Bb;^�� �L2&������ENѸA}U�`TI��[4�G1�SgXwۅ^+�ҀVfX55��#Wg��N�w�F��i�C}�᫉��h"�!�B�w}�� ��r0W��9/��!��ܼ'�|#��ZHt�p�7���T�v|w@z���	�R��<�0q��\�ci]dIx��x�Ļ�ƵP1Y!�;��R�&J�f�/-m�� �/�%'�/q��γ�F�@FK�P�$�Z��nv{��\�I��씱��K�!����AF�������?�]\u�G*ѧÿ�D����C��fW��FR�d1�	�p�UQ�@�գ�]dR:&�π�13�[�ըU�t�4�n@��%q!=������%ĥ�%��r�!�38���5�Uj�;��]-*f=eЂ^y�ӣ����n�`<��f��"���n2l���h��^��w��qY�͕��Sͦ}�p�S���|IB����ں�p��ŨV:LdՌ��F8�Aj����t��7Y\����=�8�e�%�ƽ̺�L��'FMv�g���ܿ���c��,��W�I�� �Ѐ,�\ĎJ#Ν���"��e�:���"\�8�~�-~�-ݑ��� �1��+a����p�����nG�5u��Le�>�� _��#>�0��U*�#g�٠�o��p �l(�:��

�S��bo��E�=��g�Շ�NͰ����CX@�`3@�HL���p�Ɖ�>\v�C.�!I��Ɵ�8��y[Ou��jai��a��;:�޿��`�#o���{���	�O��QP4������~[嵽��� �*�EA��O��yI;��_S�Z�a�f�~Ǆ����!�%�+��8p�ϊ�@�Ƀ+�y�i���a@�|�N̒	$z��"�n�N�?�U����(
���ڋ�2jX�G��Ch��]͙'@6�X�sا�5�]K����K%������.�&��pc��
�nF,��EHeY��Ż��ҟ� �E��1�Y9<ڸ�[��*�|Y���9�P\�퀼GPC$��:`���pP-����E��<���t�}��{�^c�l�&�g�)����q:d�`���lt��c{хFi�����n�,�]�������ۗc�[P¢~�k (��o$�J�=z|��[�9ܞ`��{��!Y6"o�s<���7@�)�^��Y'�X_ߕ���W����R�l��t;n��ۇ�)Sv'��0����ˠ�)7���:�ܫ�f(�'i�U�P�W��8,�{�X׶����
R]�!�B{HL�N6�;�u�9�zGZ&t,K>�!�ɻ��^��Y����}�}�whO$
���m���>6�H_J�H�88�R��5~x��-��>��H��g�:�������Bg�j����Fi��v���W�JP5��v�2W��LP.��%��0G!L
V�F���8�*���s��"����$���7��(u��r],4�{ c���aX�4`��o#z>~ˠ�u��IgjW�p��*T��X!��Wr��o�6�-��d"{;/iH7��I���	��:�Wy���by
pؤ$��q�Z)-��nm��� (m�>�b��㈘��M�e#�52����r�r�g��ۂ+�DI.���r�Fܺ3|�狁�DhO��E6��Q�!E�+����_�ra��CC��+;�ד�}I�l�|�Zm�X�ѱ@���hʄ�rE�BH��V���*f��l�q���C�;��!(t���1?C���ĝ7A�O�opM�b�N�*�:���FO�::��\Iy%�t~gS�K�(�}l����.wKi�7/��W�����*���헆 73���c�)�_����PS�'4�~ف+䒻��LJ�&ȭ�n����0'�Ԡ�-�j�G��^���&��D@A${;Qy��f�R��S�U	`�S�Y��(�H��?�K~9w u�"��j[Ȋ5Y�b4�|�n�)�LzN�?	3BtcH�����J�_9���g��ҚY=w����͡��?�d&��$	7��Q3�  )�"Qo��������+*�4G*�f���j���[���^/`���ߎ=���� �����Z�����ɏ�U�y�k;���_8w+͢c1��5�o��6�V���ӊ�e��FqTp�䃊�Ȫ>��X����f9n�����M��9DR���V���o^�H��-����GY��I}��1p>���K��X��O�"uǃ��%�Zzu~=ln�E$�}�+�0Cm����p�0��7ȵ��Φ�T"��s�3<0d�;CI��lq �+��%/��G��{By=N!U�i�&:(�27Q�|1h�T�G�uOr����ћf��_���0�檁�d�M�Hƞ��|N�DY���p�V\Gyg��V���!;�@��,f
F���ݝ�6d� D�O�t�\It����6y|�'V��,:���aL�Ѷ�i��4�Q�D�]����@~}t^���E>m�]�@�p�'�J�U�^�~,�_'�
�|9Z餜-�Y��6���2��R�>�`�f-~o|f
0f8��תK��.�`n���c�{?rf�@���(����g�CJ��q�T��`f�����L�%s8\��#��������J��'XV��p�j���H�:
hk�d�`*��T$�=��#\o�k�`���-��v
$I�@��@�Y�����k�R̽ÿ�נ_��A�7�)��ΧܛDwݖ(�{�u��VnRِ�c;��
��,F&�9k�%U_p�r�Ւ�Hc>�LQ/�g2>�.>p�Y��ٗ"�.�9��N�Np� _�q?ڶ���T�\�*Px�_�~�ԧ�)�D����_\wO\Q���JO��y��n~�ٳо��� sg�'?�̖��� �Qd����"r:8H�MqI��Pv�N0W�)�I<��YaQ�{N�&�:���8�\�ی����"'�1c��b8ce�6Ǯ�x;��k ��#I���Oί'^�k�^q���
2�
 ��6P�r}8���|*�*?\͙�o_m��/R�B��x��u�{�'�6�5�����]I�IS�9�D�ڜ�q����f�<��V5ɔ��77b��@S���<��h���3���2�܄C��g��2���U���&	e"P��72丑����s�-R�e��5��0c̵�G�_� [��`�Zajsʏ��@A�Nv��O��������y��»��<M�b;���E{Y��`����{i��`*��/�M�2�q!�8�z�"��-�N���De[r�}9�ރ-���8(ӣDO�j2�	��Q��+a	�8�?v*nE=���e�,K���w�;XD^~��b�U�'���0g6���l�Y�g��� =�ll� 9�@�~�u��/(�m�e��"�`Sw@���W��,~DQAu�
�?)�kiSD�(�b�E7&�Zh���k����αg�+D�c/$V6�h��&�Y9сF�ų�/A�i&6`�A�Ķ��_hp�a'!-U�g�2td3+�M��"������ډ����m8̗W&H��r�m�]9֟0!8<�'T2��A��z�n<��X�+@�$p��U$j�ֿQyO[�ϕ=�p�<� ��e�Yn�����O��U�BR���=*��>[���;��{Q� x%��`p&����3Y��{�XÔt�O��S ��ڮNi��btl2-T����7܄�'E8P{A�h!���o4c���x|��=�|*���ܜ��;+p?J�����[w?�6�  �dt[Y�3Vd�&��&���3���r:OIд�?}���p���Jt%�7t�ľ��8�?j!��؁�K�A��w.d���+e���}+�ǃqǹ'��S�|B4�
�,���W�|�E��O�	���c�nDQ�hǧ���~�- ���
]���7N��渃�aA��x����\2���SN3�73^�3N�L���}�����7o�t�Z`�l��Wd%�
eUFˑ=c�����>�i�񷘩I�� �/������[	��#�0��#.^Qn-N`��f{������9GH[P�#>g�6��c�ܘ��kc�΍�~��Ñ�#�L�;a�t_e$Oz��s¬�+f%�j��х�0��QG���U�NYlzwi�n ��֖b_!?����	%4���a@�t��Z�����JKdG�:z�6��h�iro��gD�C���H;*��*4�l�r���G�2���t�Լal@��P�� ����U����D(/��K��oq�R�.|j�C{�p'��=X��iq����`���=�C"dQs�����:S�?6Y���Q��6�g�?h����XZp/���������߫Me�o�K��L�>�����Q
��i>eLg�*nC�xG+�Qp�-ق�!'|2ߠVmrm�kn�#��z�m��|/Fv�MmF�P�����(���\�Mxxç�~�t9Uď���14%~vv�����]�R��N.H�>��q�Hמx�j�Rׇ�r�Y=�sfg"�<�����L�y�W �|���v����ao;������ =K�'�8Rz+ٿ�(AJ<Y����(?ܨ��į������~�]����f�V��v�\�_�	�hܑ���8=#1��]�~i���+qo��J�A� 9��t��\�`/�}�U8��56<qW*��T�H2?)c5�.iz(�t4�1[� �xvw��j�oag�c3��5�:�
3�����a��|K>��s%��i�76��I�aZZ!�[ �+\K��h!��1bv#�=�X�.�FdI�Yc��]�@V�C`�D= ����{��N�B��C�u�[���}�U�_��#�z�!�D`� �}�dڇ��7ަj��C&��P�$�s�򅏏y���fU3���J�y<\����cͭѢ�b���R �$�Z{�U��n�Yb�pI����!�2O��_�C%t?j����[��3��eCuM�<ɮhUoF�rL�k���ŉ\�eԕ��,Bٚ�Xv�~�e�f�&l��I@i�N�g�������6�X|0�r�J�Zy �I�e��������j���L�C�P����
#��"��ѽ@��|�4���
��$v��+�!\���JX-G,<M�R�1�n&{�M�B�/�B�:�:�ǫ��)���m=�}��86迖V��&1
)O�T�KAu	��M�qWȑ�Wx�PE`r��rސ�S���9�q��LC�� l��%\�PG{��uy����.����$9��<�5l[���`%��҈�S�x
𧔸͇�o�M���=2��N_���&�Ă�2"�b�� �;�;)|B��T�D��;��{d�D��rϽ�*��D��̎>���	4ޘ�
-4I�:GF�X2 ThK����t��@!�VG�}��ћԘ�/<��c���jl�'�|5X_��S�n�Yw���.Ӿ��ju*�|�Eބ�z�Z&���0/L3����qVo�BM�Rʑ��t�_�zL���Anɩ�6N1.�9���JO�S8�8Q�F�rb��/�ZN�2s�'I��Y7�=(��16d.��� ۋ�n����F�:Jh���s��fp�pRZ����u�4�W쬳���F¥�w�>56� �_yS����[��Gf��e��v���^�,1����� I��[hӮ�J�9�*RВ���]}��I��y��W�>���wU�i̘(�B�����<&�h���5'ޕFNK�j���R��$ś���m�aWi� I��P>y I&-+���b~Gu�諮��q���Ji<��G'%���6�J֊ϓ�wھΣ=Ի<|S7`k!�JZ�_R��ye�������t`�l��6˿]��T���e�=Wu��>Q�9`����1ƃ�Y���zo^���gx��Ɩ"��c������庺�u�A*_XM��7;$� ��]�@��שg�J��m݈H0��x bEa��hf�[��_ÎXt�<�Nk��=߫x|%>�v~�W�T�Rئ��@)�+lw	4&��P��RVV�'�ĽZ"�����t����������r�@2�"��.1�_���>O�m��P�� +�f	��~x��a�H�:��݃� ��bW��k�����O}##���� ,�_A�_�5�V�W��e:UeO1D����aG\��Z��\u��K�mQ��kdr�F�?��kᾠ��\΁^�ˊOIt4��o�����\���<�������(��~����.h5wu?�@�SI�l�L~��BkZ�X�T��?W'�^���JW��q)��ĺM��ۑ&�T��n∵���z�Y��|�?�X�M�M�Yp'���U�^����M��ժ��4��>A0��'􈚺�P�T9�+k!���
Xv���ArU?�Y��]�`��+�5t\����E�#L�#��w���)�`c�+�!�j2sm�5�h�>���(�(�RC�%,�nZ"Q.L�����!�^����E~�??Bn�����ļW�6D��|�+X��7	�E�T���KT�5O��!~�����⚨:7H�1<��map���+-���K$(�wmI!J��0G42m�,0�c�����n��㟛����r�%_�T�:�b�/9��d~�z��0��̡ޡ�/6n���6�>V�v�*�ԙ�A�(-����z��Z�V)^j�,� a,�p�fS>�)h@���}����ݼe�+v���^�O����P���n+;�01�ǆAfs5W�4=��N�e�Bm��a��IR.0!O%�=�v�fC>�����0u�u0��%�߸��n�z+5w�[uĪ���G��6< ���Ђ���|u�m%�SR��{h�ˏ@.}����Bl��5}p����)+\{M�)<�/[��q��lz�S2�䘴>��`�`4�y���λ=w15��U�j�>�n�D��6�v�yW��[qA/L{����X5%�S����ћ�i^xX��@�����,vs�B�t�ի�ͽXɬ��먝f��\$�m�?Hb�Q������*pW���ßOE��Z���.֒ՉHK�y�%�6�x} ��ld^��K�%�.�c	W���_g"W��o�bV����X����#��7*Tۧ~cN��ޝ�9��w|��ِh?@��ٿ���GGs(��8,�CݗwB��ɰ�*0��e&^z�.�@q"�n�U�?up�DK����/�k�+������|lOj���:M��.��гƷ���~��U5.<~_�~�5������voh%s�K�cıGC!7�c�Ï������������� g/R��_ELG�eY#(ta�r��!�G\2Ip�e���g ?�D��e�����[���a�K�?M��O�ed�"@���9�0�	�qM�(2K[ӱE��]�szg�$�� B��ȵ�rI&�l����I�VF,'86�%7@�N�̼�#�������t�@�O� ���Mۗ��K����v�Q'�/cv�"��Uy�\+`B�헾�e����TcQj�T|�_��	"̺��Y�ܾ���q�&ro ��r�͋4�����9����l�B��4]��$N�]-'M��,�x!�:#�ե�kB)h�e@�g!�u'p�
�ȗY�5�,NXK�oǖ?� 
Ѝ8�`EK�O6W���x���b*if�)D��{��B�L�$���Ӎ<�.�e��fP�^�e���J<�r��Λ`��ò�G�m���O�Č�n�K{��r��MH�B��9�i%w��r��x}��h�����,[ &����V��g�c��b�#�OB;�|�(�؊��rFH)�pk�Pb,`f���3��\n//��_ҫ�wӰ�*�)~n� ���u�w[�/���4�3�qeD�z�t�%�V��8K�ͮ��ŢX����L|e�	2J�+��˨R	�&%���ףo2�hL1 ���Cs��T���5v�������
MS��w_O|O9Q��́�
F6�Y�E�$;�m���5�"xk{n~z9��6��b�'G�=��&�o�����04�A���H�^�lpU#@T{���_3
d��=��j��	aġ�l���=���S�v�I����ӳ�8:�5�p�;n������V�/�X�t�b�3���!n��w���Y3S�u����v��sB{ͩ(7�����0����u�����P����O�dP��r��Do�P�`��N�:�y�7�J����V�^�ڄ/n�`y���b�x���pƎρ�Gg�<�e��O}��b�^� �t�^��j�,�ee�ι�Q��f�,��թ�|!��S�!�3)��C4)}R�W�<q�׌=��.�O�c<ު�Ƴ���Ù��D�~E���K>Og�Q3�t�hՎ�L�������m�i+�:oS/������tĵ�T�2]���5w�+Fo�eD�z�۵OK���Z@|($��,��Q߂�"{D�g������F�.�M?�w������hl [v�b�w��*��*A�gyw�ηr�*7�A� ��b����:����6�dDNP=G�Tԗ�'8��S�"���qX.)ѧ��+VzΏT�Zv{X�=��ZX�8%��>b���=���������ث<-����[�r��7}+��a �v��yG�*^2ri^@��h�̧��c�P����43���|�T�}��T�nEIh	�������ݛ\�Vps��2�GFER�ۅ{v��o�Ͷ�>�9
2�L�;1%d, U7�5�A�D��s��:?�Ԟ+H����н<�;����m`������'P���o�ּV���
݃�q,�q�'�[!
��C7���)�y�QPƃ�O]����,�XT{�[#�Z�b5���*����z����2i�Ѻ�V5��Q5��a&��.e�C�����
a��C��~C�ux-��x��IccVo��i���b�l���Mm�[��,��X�vx�W?K��/�X���c�X��2��̻wn��J(��ߌ�4�C%�Cw�f�T_�s�1��lUC�����E�]����ɩ��+�p!���{I] h@<:��xy��z�m�2I��	��UG����U[B��@�?x%g�KJ_� �*uasG��#���������Jgtr&|��_ո���hXZ��Ј��V�����n�����W=����o��V09���UdYlv�9L���+S_�R*�7���e���`@[�|[Ӹ�_�
1�� ��LD<߇��t��s'�b�������u���W�^:�S_�,i؀�zE��(�5@Ub:a{/��'E2�E��=.�2f;�&��:���)�:���:|�Q$T��Г�Ȯ=��w�T�7y_�o_+*/�� 1_�bu�x���ߩ�v����u��maO���\Y� ���O�Ϊ03v����<c�ۊ����x>�j�Qڹ�����M����,Q~��L�툓Z��
H�(2>��$�2T�4R��r���5\=3~��MX@�H���U!���\Q�7:-6[�.f��`Wc��Pj�&�b��4�M�@2}Y�s��I�	_����H̍ V�V�ɚv���Y$8���m�kc�>sy:`ɜ�F��%��|��7����I����
�o,ĸJ!y5��K�೻ .��u��@�R*��+Hg����[�Ѱ�g4�hfO�]�}���,>FE-����i�LE��1��=;!~
:��ٖ ��-��K��B���M=p��yrr�܀Ϳdvx��֋(��-)�D��|��i��q�Tr>& �V^.�^�k����y��V�S�#�ݹ���d?ތ4/�kU�4@�1���td����;�����Ďx�W;Ą2~�=�����s�Q�{k�8�_21�`E��\�쮯3u��0�:�3�;jd�#m�U�v8E��� �9t�%���V�K��A�3{q��M�2��y�$��*�vm��9���B���f�E������/Rhr��'^i��gN��~fJ�j�\���j�y�3$ʔ������P[��|�C]��H�������ԟ	7�A-� I�D�1/S<?��@�|� +g�C�g��4�f&�\�/g}�l|ou�*�ND��/��+�2��K�3{YX��'A�X/3����8�aӴH���k<!Ă٦���լ��.�"��M�.�Ȏ��G|�W\i�B�KN�Z����T���a��7��,��R�wa���+��.���L�)�\4L��J�i4]�ᗛ� 3:���/,&v��D�d�?]�[�=!�j!���ayb:�PL�;´�i��!�����#w�ao<�up����E�OqR�K�=�,P(_pE4�ց[�Tb)���n�a���C���D-mm��O��d�CK�k��e�-��Ѯ1J*qfyB4G�9��O*���3Wtj�jJTg�c���\H���_�,���Ƽ1�C��k�ψF�J@*��+������ V���_g��J������{�@CJF��jX��/�m�6.<���	-+z�F�:��tK(�1�t�{����2����ޛ�a턼�}(<I���dY+R`��їi_1<g됌�4�
�D�y�h�8q���DQxק4����`*i酱��©�b���ܡ+�V��=�O1�Bo ���.tM�=�=V�Sd���{����[3x�2�-�W\,�]�jUą� �qZJko݇��|1ޤ}�?$h�*�RT2w�+�{�]:-�n����v�"���s�U,��t����ѐ�@��R)���z�]qP$�G���B�҃GNm+~���NWs_``CUB�Īi���؁=z(�k��z�9�}f��L�5{���XK�X?���#��P����D��>B]%Z>����q�^��O�,c&�ǳ%��-~o/G&�V��+�G�d+��BQR��o��b�N(�K�i���а���Wȷ%�a�]�^oϜT/��2Rl�sU��h�"%ճ�Q����s�.ʮT�Ԫ;�q���q���д���>1/6��H���Qn��"j��������I���8�x�)uAد5D=��@�X\,!w�G�I_ ��H�{lP�8���fG��m=��jH/�LAG��f��{sA80Y@�R��:@j��Ӛ�߼�{�ڒ�K�)�U�\-�b\�!�4x��3�᨝��y�ф0z�a�A��I��#&^[~ �R0Lh�|n�&�7% {;`�����+:!�����I;��� ��#n 6N}t�<W��={NP�/!�LAM�:B �h��6�%�D�u�\�NUՕ�����Q����
~�-�)�+����YH�$	�lߌ��d��h�"!�jd��",�)�f��w�%�Z���,r�h��wk>�h�})��>�RK)&!J�e��.��v-���\\��;��>�P��B|,�&Q�Ŷo����s�\�ϻ�A�w�r��q�o<�gȥ[J+�{.ɜ�~K#���ьowW~�����98:{i�b�.G���)K�ֺ� 4��Cd^A�x2M�/k������UlBt�<ɸ �< W��Qp�~ȓ��+e���*�%=����7�m���o���C��%-�a�U��WZ��\�i�D$��PI�a>H��G�wB��@�V��������(ط�nsL0}t#�R�'�{��h ��S�M��2�MB�t|��.�E}D�,~�����8�1��2$�l���FOr��o�Y��<]��K�n�K���ׯ�Su���ޕJ�]NB�V��^��8�q����#�t����G��P}��{햤����8
c�':��龎����" ���jW�$���cP:�v|w�V����˽ ��5;�5d�I�4�5���)�){���,�4�۷��쎧��;YX�Z8��b�5k�
o� y"�q���7��r9��7���[�jޛ���_z���n�≉�!C0P2=�>yX\�OW�%�����o��Q�W�S�A��X��X�)��C26Ç4�A�`�&Ƌ�K�3|���L��D��zj���SI|w<|�t�F�KG�T0/���L��&M���HԠ�Q����m꩸]��A*��N����%���@׉��x�n�r�$� %w?ji�	x+W]�̲ �J��47ǣا¼��
��A7��zto�����S���/�FoP�Y���A�U��X�ZV_X��(���$�@��Sq�t'�"+K� �:k-~���cd4r�X���6)���#����߹�4i:�q���K��A�f��B�����2�DK������u�㑋w=7���KQ*e��Jhr�����4H�LU�tD�v8���Ǘ�T��A�M���\*n��Z�Odn�%Y�"�{m>$�qA�Q��`e��tK�{'���&4芒��HˏQ��u'��c�5Jb��:��a��a��,�,���Zo&m�p�yQb]���\�YIj�x�4��pI<) �@5���~���5�z�I@���0̉�(�-7S��&r,��~�L�P�4*Z* ��2���x���>8�>�ys���Hg�q��� �W9t ��+|�Y*0���%z3�l:���1ߣ�Uz�AƌgU�X���W���g��R�A0��Y�rѵ�h�dE������~Yl;-��d �T��^��i�$��B��CȤ��{:�A��W&"M$咝�s�Iq�����EИ��d�/aoT�N�".��5s���2������1��p�S��q�
ыd���+��`�`�e��<~�M&���c!E��<�C������a����QSd�'}���
�6.,E��;�Z���Q��]��(o����R�m�;7�E�q�U�H������F؞H�Jk3���0��l. �[Zn����/�˜6Rb܂#E���f0~sʰq�@\E�\aҌ�n�`��L�]Vs��' 5�s�~�@�M���z�*1},0�ѫ�����<��˺Yy={�3�n9�_�$��Z`{>z���������餱~��\�h
>=,z1W�p�ƶ������](s�?e)���O9��_���<w�����n�^r�����=�w�.B Î�avZ�יG����EX�Xվ�2��ȃ$*����ev�u����;،�_2�m6���"RN�\��(�N^$�ך����al C���mt���H��`*�����3��)�'�"����[z���.�*~K�T8<��lr�n���ifL]��`O�q����;}����w�H�\����I�5���̀i����2�Sz)�j�T'�
�.�j6��Dp<��ښ�w��xI4Y�y�-$�ٶ~�k�/�7���:0�8��G9v+��L7t���T0ӯ,��
-琍&��j�JdIk����^F�[g�����s��h�k�����X�i����s�+�qU@�{@1tt?~GpJc�e�Y�Z���-��>��[�:�u�X̮���t��nu�3df�R��Z�w�Hf潿��v�fk8A��b��.+8 ��tCAQå�6�"�=s�����o`��m� �=�g����X(tG�������p%5��kk���_��5R�>�=1c"ϑt��1S'����h�q���^J��%�� �Ẕ��V�A˖�6[�ɡ_]sB��)�;jA�i�,n�>���7�U͵���]��"'$��}����`�I�wb'C`�O�i4/���W�k!�?X	��=�H�z��j:�����i�Gg���Uv	S5B�/�+ϧ6��wѻ�_�w��M&�~(��K^����6�X=��ѓ<����oa!Ei���b�V���7w�H�9N���H�Ph�*��U)�=�pTL>-8s�����u�ǿ��$��E�>{��F'�.W�R�ǹ&�`�1��U!�a"6��=��1��#�A�ӍF���U���ci��Q����czk�*l��0bL�Q�*H�c���,̼VT�H���/�cy�^*�#W��������c�`z�Z��%���b �ϮDc��6����s���k�K���[T<��-�AЎҊQ�6���6�J�=AX,���mȀ���z567��S������)�jقݝ�"�W�?�L�����4wVRe'�w�����z���X���0����n���Q���0*ۓ=��_��DFs�Q?SN�J���/����ט	y̜��v�^���~��������+�YP3U#g���^P��n.eD@�,�[P�\��ů�m0�C��Ck<IN��q������~��m,�d���*�8_"J ��Y�g�A���4�
"��o��n�ͷ����4�>��Ԁb�V���PK4����Ť���� g�ﺆdN����v���J��v��ye�&W�4�5�,����=�;wl.�i6���m��'ظQj��!w�MH���u��:~��!a)�Ȕ3���af�R�Ƭ��s��@�*5�tw�mЕba��9�_��ܾ�c@��#�&��P*)ܔRR\Յ��T��T+!:fq�#kO���s��#���.&����{�����U-�7����G��f!�Q��R�0��c�.tِ`���9կ t���;bYqw?#��=��/ ����J�� 7��z�;��dGF�������)�Ş�lWj�±z_��q D� ���-{�b�ATm�&�[��-f�VV$�b{K�(�!�7��ڋ����{[.���:Q��nK�ھ���0����dY��nV#牘�o݂l�5s~�Xo�|*�-�=�X�Z���2F�a�p��������1�JG*X���a/�v�y���Tfl������-�o!T#{d�[��36�j�M=�!c�"�<��6�o�P3�#�m��qq+D9�����ubsL¾8.XD�A]��甦��;}�J�mS��V�(9�ǥ�D� @�HcJ��~�p�2�}���p���'�������1ȇ̮F�� 
�
�'��
:�>�u���r�n�
���g��B�\����ƞ��rc�����1U�>Ήx���z�xB	����N@�՛�%�vG}�����P?�	z&I��;��_5�x`8���_�}*RD��1}�ALpv������MYl�4h����xpj5Y����+�88�����@��� fH�L���� �q�Q�3�ҋw=�4k�.E���Xi���C�6����͎�c1���k��$�Y�����-�>��)K#�KK���9�;w"Q��~|�|,X)6�=��YEɛ���`�,كxŰQ�k��C���o�փ���+=�0�F��3u�$�ӬQ��W�܋4����őKLn��D�P8���Tp�_�cҺ�������1��D�th�2�iߖΨ�H)j!/��uݪ��dѯ�~�\�XB�����;�yMss��	����2I�]��^�ܜs�]�Y ^�[f��M�J(�5�c���L���-QӃ�1�.��j֡�lp6��g�
�J��m䎼%l����>4���vͪ���T��`?�~E�w���~<��Y LX^�l]��V�O�TB���rX��C�7Dv��q��X$�w��.����N���JB��h��	��]j����a�fz��~�Hk���`#�>�D���� ����h�>�cA�ָ<�����  ��ꖵ�u���S�,]״~���K"���b���[�j0q틟1�\�l���:���P+�1�{~x�J���QpD�������eG]��'��]�A��<���qf�3� ����d����)ǅ�r�A��FQX���VS��'��J���e9D� �肜|�J�`z-����Lb"�,��q�r���fN�L�X���0Txc4������5y�q���;��r�"�&2�'+�*�T_*��ɇ��窕��O�q�Nӱ�B��9���Q`�(Ӹ1�8͂�4��N�X����!=Y��� ]�t�@�N�*:X�l�D%&��g��d�/��j�W4����C�������X�i�<���gV?g�<��W����0o@�Eߞ�3*��}�/��ʳ��4^��#'�(��<k�嚐/����$�"t�ue�;�\���d�w�]aI �\C�e���}w��4�z����k�L�b�U���N��=Ė�`RX�J�������E8�F�9��D�O�τ�n;}t�����r��yP�;�@&�t-�Mi(�z� ҬA��ݔV��x@ƃ'۴������v���GCH�S�aF�E����-��֯yȺE>��E�)� ����T�;]��"g� ���Cf� 8<J�O<hE���{-���H6��ti�,)��	�
���$�߱�[v�[�a�$��q;��h|"��/�ݍ��ԃL�>G�{��bסn}�;��K�"[�ӄH!�隷�.��&��ƿ���q/����C�V��9#�$������6��I{�4�g�Z��<\���(������� U/ӭ	5wӺ]�<~�ɪ]h���!�#ӌP����y�W�(W[��2|����t��0����F"��l���D4�r�ϕ���GU�[� �/�4�{��C�ӻ��k�Bz���|#}*�	����l�[j���|�<��4�N�i����@E=�{� 4vS)wY�C��inPt�|��ʹT;��B��&��#�5ÞX��-G�r��#�j��K7A��1睨��%J|pv�e����;<{�>=9���&望��Z�C#��)F�㚜��X8N�'8C�;m�ҭ�{7�F��d���B�c.TG���� �k^���T��c�Zqo����H%�[[��w�\o?���x2?��Z����b�5t��7�ī���[�o���9�s���:=oƋ��I0ζ|��̪��-�j/z��6(b�$���C:����'yp���-�ט�M�Yn����h��I���.F=]$�_Л�-]u�Bi��?�tAHT�l��pY;&iw�%�{�s~�����Q6ǰ��/0��y��z��ë�O>h�.�R�GV�w�\cCm�8ч���2�6��S� #p�	W\+Z�(]�X=v&��?JJ��'fK��v��u�"Ş$�pI����<K�ⓘ���Oi>h5�,�A�
��e�����M������'��#�.\�⩕��[Qj��گ�nVh�
$�!ׯ��0�6���M>�}K�+oR�(��\����gÿ�'aۖ%&�
r��`qd��&ʕ͕���ɭ�Dz��o}tQ��9��V���g���=���}nA�8�")ԙ	�-�6���6�������Ř��� ��}���������|�@u��H妍�ؘ��1��B�ho�z#����N���ʢ\g�̏9�=�m�$����U��_��X��.�,�ј��O��D�\P�|R�����QF=;��Ep���u�m���z/�S���.+�b�A~on���B���@C%�.`1�I�DnE��;Հ���ըw��j�.��?IaWH����TL����T1��p6�(t*Z1��&�iSQ�7.kL�ySܖ̟J�ڍt-�h?�K8���P�+<���ʱ�g���W�I�����BaN��W�]�񇉵�����DOt7��Nl�^�I_c��lV
����B�v�ͻ�#����;��J%&�Fs��;�YB����s��+a�Pj��B�֌y���Ya.Т��������7>���>X�##ݖZ�|�K�y6;��̌\��7�q�3.���7R4�K]�u�%9��h�z�E��r���N���  �����_�!�FV���n�h���X6�X�)WĶ�:9�#�R�ǡj{�]Z%��`��E�븏%�_�$�4�*<�ة����L݃�.=b�x��g�I�{,H����I0/���!�O�����D�I�f[�����Yہ��v��������̈́[+����I�o���ƀ�"��7'`�X�L��b�7�D��~�<�Vul$�Y��#�-6��ISe�M�x+$?����p��-�n�z�)�?���Gs�&����4��{d�R�1�6wٟ��'��N4�4���֪1��!<^��rG�z?��5JL$P_p�������F�f1	�
�C�G"�KŒ�U�y�ĵa��ڛr�^	��GNmF�C�^ 8��C�(���o��a�6F�'Hi�-E)�J�����ͪl�E��Ϛc����G��M�\�����|L-=P�k��߰���8�E�?
"���5h�*<��݀2�=��uS��WPYՁ�LD�א[5ĈD�ɢZ�1Վ��f8��&v�8��GͶ�nѵ��li��a�B�[Y��m2�#g(�T	���D���!��T�K��?ߟ:�ƿ��*�������|7��L�@l���=���O��]��F�{�	��z�����,���"�{���{�즻����(�f;+��X���7`? �U8Y�w勞COR��f���%EO���0h���IC�]L��DrZ�0.D�����{���/i
�Hm]���ܤ�K�&�E��(:�!����;>�uZ@�-ʂS'n���O<e�
M�� �H�u���@�}<�"CU�c�����QTr-gX��Iw�r�[�{�z!C��������Y���'"�DM(�	5����ji W�,ڈWk�"h�u�Q8ڧ��h0���׆RހHL��=<�뱚��`Gfl�%�-�/M��F;Xr��dQ
=2
g��rUbv�͏]��E�`���Kw6�Pm����Z���'�iܝř�9t�^5��n"5�.����˙�l2ۑ