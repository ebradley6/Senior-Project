��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z��4֬��9�A��;Un��Gh[�����<�#�L�-8�o����X0v�c�4��S�`U��� ik�{=�g]�C�+a
>kN}%]q�]���g��k���Y1b	 ���5��G��r>��T�CF����Yf42
!zEKǍ�>�e$n�i��F���C��T��:�/�ig�Aރ	V�j�e����@Ȋ&��<�RL.kD��JQY�q-9c��|�e5�P~+��q��ͬd�[��@�A�cB��V�4?AQC��.4�?�gI" _�{44��!�p���H*i��˘�$ǴpH?��Ym��b�H���ёcd�^��RN�;e���[��[�s��O*�`e���gE�rh>Gܹ~6F���A�9���uol{�� �)R�r��JZ4��l	e�6lC�D�T��~-�H&ְk�i��(�Ue�O=Bs�����*��jaΙ�p+��Zrܼ�-�1Q*�h������8(��z K�hR#�]��d��p�=���Zx��=!�7a)/�}z�'����w[�SG���",��#U蘐0�చu�G�[�k���a�LG���2�r��z]���7x�Ɉ��m�T� �O�L���b��9{������x�l:D�9�l�]���gh}�6\\z�G�du����I��t���1���Ȇ]U�2	9�_j�����J}�a�T�a�=�����"2�������N�Y����I�q�D�����u�����VU������S��=��HJ�1@�gj���ڈ
EXd�@%��L���D@ef"�2��82�ԅD�Q�5��"�B䗖ɨW��gBr����t&
��A�aUW��Q��Sл��:�"+N[`w6K�:pA�;�����?�.B!��
�,��?�>&(��H�g�L�DYVy�]��d�pxM�<�'�%+'��,C�(�1�����6�bd��0��F.v��'�:ݤS8�Ew�bY��*��� e�C��$��w83��e,���8BM`�U&^ig�ǎң<Vn�HJ�"6Uʑ�fJ������X�ρ�#L�-w�J�r�[�۽x��9�}�|�����h#m3>
bE�e�a�#�k@���WǷfX��/�_�\�v]���UY˦�a�W��SB,HB"+q�Vz	e�s¼��nM��>��k^�e���K}����t���عN�m�ۍr�u�	cqٓ����������U��:�&�Fo���È-�|���-��9_s�,z�$c6i����M|Ҹ��^�,��$�4�f����̢:%��9�$J�,�ְ�P����	/k�a0Y�WO�?��ğ$�|�@߽��JAeY����͒`������ᓢt{����ҀI���KƐ )�W��BW���e�G�C��W1����Pu`4H�\��`L#v7�e��3Y�`������zz�8Ni��W��F�F��^��֖d]�Y���9�Ȍ�$	Ob������_Dn��,�Xa��v��6m�m�/��y<V�WpÍD�tx�vt�ᢱ-n*�6�s_�X~il��F�Q�g��r�Ξ�r�b��$��>�Y��l"*��[��'�n@���i�,vb����V�E{�uW��%
.Ҩ~�Fk�^�H+��Z^�����{���:�o#�����@J�H��bٜO#]JM�l��Q�
La�"p��M��#�,���(2X~��q���R,!\I�H>��(3���ҹ˴TrQ6S���9�g���_QKf�=fP�"�����Y��6�T�ֺ�$��KMX{�Lz�D/�͈�#�H<I#�����Uŷ��\�'n����^&�5����#q�
J%�OcK�S�X�R<[�H����*������Ջ*r�&;5r��ݦ}}yS�[ݩ3�TN���pw [����vu��^j��-�.ZN	�~�nA�#���:DDĕ��Q7 d+2�b��_���a>':.���;�.w����_S>��]� (��S�)�:�+�|��|��L}�E�W�+!%x��%ȪZ�'�Wr�?[��[��#��;1�A�%�d��q�����>y���Ť!�L�Kl���]�Dļ�t�&lr�����y��?�������
g��Nά.
�$���Nb����v�Ӭ�M�<�J}�fTU	[;��2����Χ�q�Vz�����Pz>V
�7���^�=7nM���s��)#gӁ�ʅ��,�|R�&���3�jp؎Ո�ޛ݃1c���%R}��X{Ɏ�
�@}���{�*ި�PU5Sb�:���0��DC�0�Di~n��q$�
M{&��2/y� CZ��\���`hqO��A�Sb���e��s3���>�����V�3O�+M3����}�Zc(6��s3$aQ)qU�a>H_?hU"sݖU!\Z>��k�ߊm�5M��4���7=>��e^�Q���4n9�4y@j�{�:L߲�L��9s(%5��qĶ X��^Jj���d��^zx����G&E�@7��iQ�O�b�\ˍ�|䒗��"8P��]�-�:��G��I<�.t<�����|,�{��r���~�E%}l��~��b�
sb�G�N�y+z�1�1x��\�w8nQ#ɁwE��l��~�_.FB�hfR}�Hpt����~�'�23w���j�����|��ȵFô}$rߧVα %k�	{K��LŃI3֔y<���VnQ��W4��_�@�|co%���(z���}�bR9�"�AGH"��0�+����^-�7�ڃ��(��*tlE�%����k^��2�EH^�?�^�A���
�f�\/�[__ܧ+�D�k�J��.b=?3$f%�8B �K�^�G��b���'= �� ��OF� �}j�3���>�@
f��Y��OQ��K��lf~��w�9��H@��$�Y�9LV^7sZf�o��'KS��*������?P�v�KXLZ�"�^�'��#j�w�i��}k$��Rv%9�QR�O�Wu������݅/�כ-jk����7�쎹F�GR�k%.����PT9� �h�}��-�l!�]�e���̺�x��+]_~�>���44J��J"t���w5؄����E�f�ѳ.��Ԣ����MC+AUZ�gw{uD�a��O0�sC7sp0�OP�)�����M$�mDǎ0��t�o-��?bTZ���h8G���^oㄥc2m3%R�&ðM�Ǘ����q`��ԟ�>W@�������fX7��eo�h�T_�<����f��[�"�S��z�����D������jvg�	�Cn��<w9�<b0��Rxr\p�2�y:m�leA��RaS��Ƥ��+� 3;��b�E��Ϣ6���+?�5u�=����{H���f�x��q�.G��͝t�$�t;�_�+�1!R���l9\�L�Z��Tw��n(�S��z��������Al4ۍ�V@��E���.�Рy;����@B�xog��9��W�}S��[��35�<e̦F 4���g\�,.�J��N]�\>�N�c<w؂���ST�w;�X
�!0>��ݕ���D��Ks�n��Oek���D�W��\�9\^.w_+�_���yO�!�M��^R��Q_3/ѵT�o}BL�?f��m�m�?��%j��t���x�y-����J��c
��"5V���ϵz�z�s��oCΔ�ì�!̰��9��M5�_��D�2�,��!CF�MEv��jD�~�M��ɽ�@�;�@)�aH�d�2+o�$����P<t%��H*5g��u�z���~��L��9c��}��'4RI��j>**&U�Yn����O���d;���'��X�Lq�oz�ڭL=6��N8�|6��6o$�E��>Թ� �������BTnu�D��gcz��S_!��Y�2�M6��@��w_[%���qhJb|J�k\��J�w�W���Ń0g�'"-��,-��6_����C�k®Of����T ^�����:_���
fS��������v�,n��$������?� �|�@9#闇�!'1�
���	雛�=9���eN�C嘍�C|փrr^�<P����o"eϋb\n�=}�5(�u2�Q滺��f@��}A�T�0E�2%{�5d�7�@��Fa�,�U��������$�
�:=�Q	��2FhNƉM6��)97*�FCZ�l �PȌ���~�ASA"��ֽr רf#$��ؔ_*�yv���A:䣴!��V�š0����1!{�� >f�w!b�˹LR��3���c��S	_4:�_G(����H$����s���xA�nu���B� &�|�r�D<ep��wd���Éhvl|���P��<q&K�4���f~��]�k�2+����M;��U�4��v�L�VAW�m�V�J���lFj�\K�2�1�n�u���Fd�p�h�R`��KR�Dm�[u���</+�*��Y��j���4�>8�i?�NU��f-A.Ki"w��c������x5A��`��~ �q"����6��R���`�Jl��70���Լ�{�j2�ݾ���;�zg���W��G�:5VC�3(����,�OPA,~�xjj<��1��-��v$��������z�K	��}���7o��o���b���q�G�T��y�bD�_�U�.�yi����a�[7_�OjHGL�=g�ۑ��[��t��4�*ID	������d��nwaI9\4%H�<��fcCH���"�f����&?��]�-��H��t��.����^��[
�K�%A�V��_h�5�����y�P�r~J���;xT�-�u�`��?o���Ë�[9G8��fw׍l����6�˼��',5¸�"����u�_ְ(΂�{���6��[��sz��O��2M6|	DO��
�OɌ��Fu�\�A�7s�H��B\;�-��WjXo���74kU�~�Ƣ��%����}���c�aL[(lf@ֈ8b�fTp�l�;��[V���X�P�hx�pPp�;l�:��(��'�]�w�ב�W���f�(:-���e}7dT��q���`�B�3�̅��Dn�xV/:A@��m%Q|#��D�`������Q){�g[��#=1=<�������K�C�4S>-Č7Ϸ�DN���j~z�%�dڐ���޷��e�˂�&Ë�U��_����6�S�!=䵳F	�Q����:�6P��B��^-����R}��;�7}�מ4�9`�<B:~w�J�����v:����-����ʌ3g�^D�}�3A:M49wQV����Pm'�y����؉�v��\3I��v��|�>;�mH�5��ftr��/��?ii���O��m8�|�J۷4{tEqX�m�pZ����$�Z�.�ӟz��S�=ӭ���͙�
[`����aps�r�V�<� A�mu@���ι;�f�L�� Q�����2�f������R?i���v	�8����=��Cr^(9�H-��K�5���44��|i� �<#í��!I&кK4X��e,[xJ�|.�mz�*\�J�?u>={�,?�u��q��#p��O�'Ǆ���YHdņ���q4�;�>Gh�y��lv<y$�wq2�3�_Ҭ��q�A����)��V}�ͻ���r�T��!���f1fL �)4ve#D�zN�qT�,T�G�D�'��z��]uJ�J~��<
����b��4߲��i����$���`M-x�KslX����{�O�Q�L�&��)n�R��P�X�i��ޣb�U�\�C�"נ��ZK�U1��{��8DA]��`�aB8z���q���=�`�9F�^���o���2�- ����z4|ouv� 5�	Ѐ���l�&�$@�9vI>M[�5��F�2�r_wU}�=�
��kޥdo-���i3U{.Q�(�ŋoŕ��C�d�����Jv�\-w(�Zd]#�!��gj��%&��-���
��� ��mΞE�Z�Ί�7��HXuro#���ȡ�q���Q�T���3+嵱3��Ā&Z '����)ȱ�vn��A�Щ4��s���|L��z�wʕdF�Z½ۊɍ�|}�L�Sݠ�qw+�XL]��HSM7h��Sx{�X��pՖ4,.	��3_j��m^�i�rP
�.�	�3-(�ǳo������w�Hk�3uC D��b�DV�J�����S�VWY��o=��7(0Q����[k�VR%�;I�w�����19�&�̠��~{�+����5X��d�EX/��q�������'�-uV�w���m�H�4�P��<�ź��B;��lKg>�:�1O�vk�l�t��Z%9�E��C�f�$�4凕�2)p�6�M��-@�h0���M�
�pb���d����b��4����ɕ��J���O�󂊞�Z�̝��e�,�ׂ�\�Iq�����dؿ0�9��	�ڮ-��h���c���v�����K�q�뒡��{AR"��2�p%���D��	���v4׼f�b��T8I����uP"�q	�?��Ø�C�>���������1G��7���GZq^��W��p�(���\�f��:�y����b�k�����*$5������R�&�l��Qɹ�����C��<Ћ�R,(.L��v�+�	�~��3����B4��� �>��*7!�)�p݉f�4�=E�Ҧ��T/]���N
.����ê����$�Vx"�kC���(D�뼍��u��r���wc������;^���Py���a("�\IY叟G�h�@�w1$��I�	�e]�NP��r��~������5��1�	b�OP�Tf*�{`��523��I=�Z�R��7�l;ІO7pw#[U��7�-g�/�>�g6�ù� �Ϧ#;_��k��8I���p�1��j���9��O�ך[��ᐾ]��-�E~���'�1�'��ɠ��(�OE�B������P����V�����YD�Ek������,l������z<�x��G"	ղ	��������jJFً��11���
Ň4C�8��
 ��J{B:v�E�ڪр�?k��9�gh����4��0�8v܄HlP�ު�jm�dE��N��R �U|�҂ɦ{�jj}�D"��R��PE,���KW�F(=�]ys��`k�"E���M����������w�>X�gU�|^�3�-2��t,
������
���鷑��;`G���yŇ���γ��FU[Bv�Z&��h��`���_�`j��^q�FY���,�S�
%�8j���)�֓�`'�v*ɩ�`ָo��E�+8�W[m�����t��3��lL���7�8�8h!@�G� ��j�dh��8`���k4����=�%]ޓlq��Ė��
��-c�\�l��r�u�UJ�\���9V)9�����v�8L��$�/���
Hۓ�d�q]��/�)vޚ �z~G`�A8��E ���%�.�86a��q��6�Dv��e(�T��=n{S�_����Zo%��/�B�ҹOQ��W�i�$�x���y�π�l5[>&��U�`�Aߞ�՝�8,�"�!�J�r�hl�o������'*�d���B���7t��v+3�z��ްt��
�C�!|���]_����^�Д�A;'h�[y�		(B�NI��1���[��iJl�r.��q|P�p�	�/�>Ӳ��B�d4o��Q���;ɞ����p�/?9wm���R�!ϟ��������tБ�j
���<߬� G��ߕ޸p���Ϟ����Yt]���m|�>��{��7����8��K�%{������'��)�@	�;��a!p�ǆ�Q�:/"C�!���j%�Aְ�� ��[�Uj|C��ԩ$�ϛ�	cL��7u��Y�gk���sТl�D�*��7�m�f�"�g���L��>�����a����&\�\�#������ɹ���*z14{�4e?�L�I-<�dI���'f��O�hrY�<�M�C�<LHȗY�V�]�{�)Mү���,5"4�j�5��Xw��)�Z�xͩ��%y������6Y�m��T��*��U��-���>1Y�Vw,h���9������M0o��-!/�ݨߎ^�XK���n���(��-�w���g�0s��+����۪��h6�:>�UB�Oֶ����U�i�nIY��\�$���z�;�Tq�O��-_""����T�G��=l|c��s�N4�b����-�|&�垛�un?�w�c̀>y7��;��ǃ� `L�S𗁖B&�@G];e�ƹBٗ�k�ɲZ⧟-M�gw���D">�r7��q���
W����JIn�ߗ���c>�붮a�~�˨.ޅ���d��m��۞Q���Z��cY�&����	x�@\I�D�󵽙���3��o��AR��&d��[:�cN�P!�`M��Q��������_�7�gv���@�3#]�#v�����8^cհ�_*)����Ok~��o�!X�a����A�D�c+���������4C��@���9"�� G/K���4>0�~J��T�kL�<�ɰ��s���x��������~z�vTP~�/��PW���h֢�2cH%-zS{D��0���\����ryD:bR�|��#�`Zɖ�F��m��K�nB�b����y{^֪�O���~!�?�D�r
j����`���m�#<Z֬�+t��˲R�:4�_��x�Gr1����@mf��6�0�δk�.�d��wB�K]qp�!��c�7
@m:щSfs.�?-&|k��u��E�(�E�p���?n�T��MC���;�{%m-UefZ&[k�12�H�=��uK1,�^���	�{|��;?�l��ueHl�����]��n];�:�R���M��C�g�QV����4G��lsu�&������]�|;�C��np��N�V�$~q�Y&�����hNbj��xOv���?|���n���߷��F�r��O٧mp���V`.#n�]�v�+�P� ���O*Ȯ�d�4=��A]j��Ģ.I,��F��hӶ��@ޖ�J�����i�Q��q�t��x��Nę^��Ce(-y����#��lyu�?���w	���T���Lq���[B ��C �+8�%/m�9*l����:$%��'��zQ����+�nI��H�I��Q�`�[-ƚ��3;.$yv�}�ƴh�~�DI�κ ;(6�5C2Z�~J��Xҝe�cc:�����)a�4ɼ�4A��b��VY�5�_�Jx�n%��M�f��u]<�KbQ�O���iO�:sKZ����1:�
��Um.��Wf�L�s�ϼe"�� 35W��I��b5.^���J���B��!��mն7��8��ah\���q�h�����-,��(�>�������1���of����l� �ҩ�Y��T���v@y-�մC��Yi0_�����Ǽ�4�#�S#��b\���`��-�y��S���7,l8�����l�`�j�����l�ʶ:�jkwh�(�Q@��˲Ǩ��&�0=R�ߘɷ�6w14ԉ��}<.�Τ���ˢ�ߖ�61�F�^-���D�K_+,�~���tB�d1v��9���Y3�����y[�P 2?N�N
�uOGG󵻡|�~>ً�I�����h�IH=��Oo� Z~xLqo)��9���$q�B��rW6=�̆���bQ�D>��%��aB�X�1�/6��nCs�������ا�E+�%։c�)e��7�pւ��*�����%i�e�ǂ��܋Q�m���o7�P z��6���0Q)��l�����%z���/N�$^0�Ý1�B�&7�/& N�1�d@r8vw�P2V�Ge�͋�;��03;�%b#�ݻ����!�~Ơ_����y�."�/�a~jHZ�T��7L��7���OB@;n䅅L�:�Y���4_�4���1F?Dh@U\�[P�V���^d1�]�ܴ���}���Or]V��J�\)GdG��㹱'!�t���z�����!�^e���in���"�#Z7�MB���V��;��CJ�0KA8[�@��C&��/���W������,� ��Y��ټ�E�T�9 NmY,�(��P�(��l��������&���Z��!�:�r���,�m��WM�ӭ�@��?�-��S����q�v^A�Z	�M��+�ԯa�]�,���\ik�/���{o�k�]A.Eݽ�_xaYwD�N|n0GS�+�%�/�P~�:{��U2��rxB�[�\ ���U���ǽ	+e������d"6&�=^?i]�	�x	8�� �(Ս�&��Xa'���x�e��b������M�o=z�%�GX��诼��DK#����3��Vm�P�n�욭NQؖ��9����n�QQ�,CİB(�8��l����2�U�N"������_���W�ӆg֥�kR�p΄����RS"\N.Z�H����:h��x��˒�-#,_�er���	
,����ؗN�G?�L퇦�}�^[�Y����7��|����p�eU�3o��Ԁ��$C����xn�`P�W�������GDH��V�_�0�L�s��C��RZ&�(���_�o�lOA{�B��#��q��F��d��ӹ��� �1���-�8�2��0��b�pn�4�}>k�yv&.nTa,����44P�0d��(M�DR-@'~ů����JT��q����yu� U�x[�j�\)N$��R�!h�w]>�z%�<۰~��<��T�(m�Q��~y��&CQF���?_?�T��A5g�+ՈE���o�j���¨i⩖=>���ٲ���n>Y7Xfa儞��s)K�Ӂ�x�J������Za�֥1�+�uG��o6�����\�Y��/(������vs�qA����V"��l(T�'DlHq�갘Fv�zT��UQ�����Y��PZ�v]
7�t�m2HW"~ܚ�X���A���L7�=�wZ�ir�K� !����4��,|��:ED��d
J�{�H���H��%��j��Z��T�f]����,ِ��9"��Ђ �$*�Y��������/�i�O��k}��B�h����'�"z�,�2$����7�1(;�Ւ!��)�7{��*�A�EIҺ�<�ɏ��8W$���И�&��ڇrh�c��4��y/JV,6�~/�%j�pĈp $�k�_~�W�$�Dˇ_q��@\!�-�	:�FK\�Qƀ�iޘ\��:�y�E���/�z�� ��d�U���b=m��PfI"f�s�x��1�9z>C
' k�Y�nF&x}��@*UY#�]�&C �@�Q*&m��Qd/f��E�r��tb拹�.��.���l��N2�F��%d���4~���s/�Ŕ�)��}#��芃��P�FWH>l$9���m z���-�{���N�_��A�y�Ep��m'�~P�Ш+&<��BY�����s�I���A[s*G��f+��n����Og�9�� �:���r��;RP�<�]�7g�y(,r�	\܌Ũ��2o%c֜U<p*�;s1i�*j��ƕ���<>`S��@�b��\b�gZ�Gh�B��i�A�.6V.]����Z ܾ��ݰ��V_�~�<x@]f3ou�b�UO�����֝�+G�ٗN ���g�5�9�>���9���j[�5��?!aDEÇ�R��0�7j��ޡ�x��ueuNh]�Z�P=K�!6��fpN��%`���� �(�Cĥ�Gwr�-��@�|�W�����1�q"����v���2�Ķ(���G��<��X�	P��cz��h�yNY�9N�S���v��Y��{�<����G �g>�K�&�l�W�8#��tM[���Df̾�fk� �Ly�N�Ҽb*͏�<U_c����&��������5s*ԁ�{͚�g�p�l(.��zo�������d���}|�j$�����2ɘ���s����6c��Ȩ�@��˒�Z1��$�N���d����[��b��W���Sy������ɽ��˫�����穑!C^� �-wsF]	pY�(���y�鄖�d{t?�B����������uۘ;ȵ�oqWT�#�%��J���M�V��F�Um�2u������o��5{�(y����*�y���=���>�����n���9_���.�A�4�b��PZ�Zc~�ã��'G:����ʴ�tb�e&Z8�k��3$a,8E99�6��8�@ ��h?�õq�l`�X�/�hcp�dd�yaOF`���v�`���#���t4�6CZ�l�|[>>Z3�4p
��4�ձ�cA��!"tt�2��#�[;_xy|D����^������I�M�55�� ��u���d���+�t4���S��%�t	�Ϟ3UPӢ���T������9pY|��/��U���O�P�R��Q�gH"K<7Ȍ�)j����vZ��uÏ�<�O�9�	*��7���"������~[�*t(NH!Cw��k�-�����c�d(aHL�lGdAA��:�)�PG��.o�T��,�]���բQ �H����]�e�1a��7 �'�|~3<�խ�jH�r|T�MGSqj��XU��@�)C�Ø7Y�k��Q�)���,�9��޶FD�Mc}����.O�?���Io�0a�������������=��dw��6whQ�ff�5¿�������N���뒉�y�U�b?�?j��}z�m��<�w���߅�(Qj��Y��i�D�3��3�7N�"p���A�+o�2IX�y�K]�T��Zx�UAQ]��ܘ�Nv�`�>e7k�]WnN638�u 6/6؇j�^s�y%��{@���L�NT���O�K������ڔ��~G2��g�Y��k�G��\�}�1,�����+Y��Pt�!(NC�k���削�����z�D�q9>Wh�P~8�LqT/|��Y���D����^\Os:	������M�;����j0
pzޕ�H�V�-pї�{�t����
S>:��YI���9X����,T�����a&����P�ߛ?o(܋�t��RI��lcyoJ<I�GT1.ʅ�:-ey�	~9%n�ڵ�E�9cl�"��s�����so�J�����L�
HMe�*V���s�UI-hs\�\L�!��?-��� �bV�S�ǁ��,���݄+�Bިڀ��D)�|�,e0F���4d��[�𭐪>u|θu����d��Za���������$;:�G��-���6�b4�&(P0n&�z.WR��A}j����CT�m���uS��%
�a�Т��D�rTm�Q}��ۡڐ�XT�`V�J�uRj2�ݦB\�tKt����dT��s��p.;�!��W����M�l���!��bS�Y�k��^��7��΢u?:�Uի����"�T��o�<>��q�:�ݥ�G�Ֆ7bdʄ3�A��`����!�Ug�'J�r"�_f�F�ER��~@�ʠ�v;Hv[�("�cq�͠E|=JH��aͰzF�He����hD�g~9(]�2�������f|�{������ m�q� x|�)�+a���%]�,-��C�7�"F٬)�����!��9���[Fz� .��?�̭9+щ�RsF@�z�$�\�ȝKR�2u���c889�y(V��$N�݆���B�.:���ɱh�������evס[�ֿ��R�r,nx�����u�5��O6B�I�g���������+��v����@�-n�c�6�.�W��y#z������(�sŔdPۊe�������Y�kms��:i��tpܳt_�}<�L�����f4p����x��?c4L)2B\a2�$�?v$A���F���ۅ�Ŭ��s��Щi�E}����^f�n��9�f|��U |<����/�P���S�Z��7�a�>�i����y7�w,�V)������gd��
?IR��ՏxZQO�8�J�����߁y)�^�+��ñV]��'Y�k�ƪ;���Z�#Nh���M(�s�ψ8�冴`j5j��i��x?���O�u�Q�f�Tvt�pgɚ�\}��n��!z�"X����d�d<�8 ��VU�����;w�o&��l�u�Q��aJo~+q�\i�U��6c�)�ꜭa��#tY�j�u�����q��)�M�i�]Zr��Ӥ��ev�gr��xы��ܛO�b����DL3�ڻ(��n��V�/�jFR5�[Ө<Q���z{R=�=�9,d��+%������Z�����{	j����i�����
�%��f~m2�����D��<4�Yq��®�;�
����7>ΰx	��Հ�7��u�sH u�q��U�8�̬�tAe	��G�RN7��`��4/k(?=����4��_�N����<��Ce�z�ԯ!�"�Wk�5g|$�-��������X��C��5�[��KI=#!+pO��Λ"E��YӪ����1 ֔�}SC<:�x�"��Y6S1v��S!����y�GA��;~z]�|����Ypc�nU�:1��h6��J0���$��+o�*s,N���M�o�\�����7Ǒ[�˶%�[��M]�LR�$Q�_�n��5�&-b"�]��kd!�6��,�T�^��vvH5kЬ��K@��|,�#�%Z�o�B�,�40�^���"##xaE= fu�1�s|D|�fq�/=��Z����Y�(q�𽁠��@P�)LF�+O��#<g�u��#_³ڙA�I���1:���Ob���ˮ���x��5K �מ�U�)���pst��k�m���T���/3.[As�R�|��=�c����BL���{he�<�_���/6-Kbi�* ��j��d�+��q�=e�b���!b�đ���s��y�>�z-���v(ӑ$YѮ�V� �=� �)ث)Ho�
Yc�a�S���E���Zr��Ӷ��հ�_�6�"�44\�*vJ����������`֑��RB��;M�~mnA�ֿ �ֆ���p�����\����;��!u�:��pj�kۧ�h�T$0�eqU;��?����ΐC/�;{�^,Ɉ\HG�z�������k�C�G�ޣ��N8W��zt� Di��hF[�!sYLZfދ����<�����B���3�f�5��A�E2��"�}��E�P��U|`J�L�K�<8��7���!Y�tz�JZ�#��s�Vt�?p�z����0�]���4D�J���I���������͵F,��h��3�`��^�Z��ֳl�@C����5�%F����z�FP��}!�m�I�(}h�\�{�l���J��h����&@�� }�h�NWb�yEك�[?;r&tε�Y3J,��v�둖4�8{���~�1O4-4�jS�v4Y���E C��l�m{>���u*�@�Q�8u�n0M* =�lK�w��.�ݯ/{($�:H��(d��a׀m�0�Qos9U-T�$ A����M�ㄡ��$����.�Wυ��H���PM���L��}˜W��K�P��j�ƴ�P=����=�d UAɚ��]j����� ѽ�A�
�7vP��#��y���FP�-���%����#g���O�@�ɉ��t`
`��s\=�N��L���#
&Z�2Y���y�����T70��.Ĉ�]'��i�j�3<�́|ۄ*�C�pe�;&UG�q9�M�}߈;*AIDLK�R���>�[
�z�1H�����],j�֡�h�����$j�B�~=��^/���\�1`�C�"͉�TO
~~"����֮�m���H�"L�u��J���5X�[� ��m�|f]��Oq�eQ��g[�Fz��so���_ *�2��i4�,
�?�o="GO3jhz�ڕ|�4�N�F}j��h�c��#U�5e�j����q[�U?q�%8`����?�D��'��'*{2�	-1�[�u8�m Ԓ]g���$�}��I�oZ�S�z�;��N�`7��v��-S.�5~��Zx���i~�$�� ��\ʩ~��wm��0~�WrP�?5gd�I��+��2��.�"�FO�q��y�?��k�Cm��qkLY�<��fuG�~���^;b� �0H�$��G��k7�r��%��ZlV�����P�b,�R�KrRWn��ȡ�c���>7��=s�����-�tB�������N<ʜ<s�
`e���t�O�D��z��}��Ϊ1��#����^˜�Qxޓ$��1����Ծ���i�j��(��a���g���D�`Sq`h��	���Z����2ǘ��%��?���n`㉨�U�>��I��ݵ�d�}��m&GΑ�	����۷k�����z�W;����k�T�����*�2I�& ��bm��N�q�V�o��u�#̵��!���f�{�����ͺ�T|zOI����`ڬh?��վ�~��$ ���=���)nJY�ɥY<Cwz3n��r	�� �l�6��E-a�(��8	5T�K���K�DVPTH
�>�jL��� '�o#��!�����g�
ϰD4~��Mc�E�&]"���.%�
����A�-Xxĩ<AԞ3>���L���H.i�sn-�f�o��(�jÈI�Z��,}� ��.c��!�6�)�tm�uݫٗo-�� �L��r�b�]W�����N��3M���|��xi���Jk9���+�IЛ��"lR�+��^���D	���L�fG~$dEB�y�閉H�q�KF !���^y�}7�������1`t�#�*<�(}�3':�����7��7�kb�$��s�Rm�X�	�6�58�=�i3΢3�LP�BI���F0��Jb�Y7�˚� \j8�u��[�JG�5;�n��l�b�)�&�oP�)I��#���L~�4�R����9WUbG�gZ������w�:����X�;�a���V_�lۛn|�=z
s̆�@8����_�����L��)G�Rx�6(L����'��׀x۫�0��S��MF��L����
�}���8-�Q�y���
�
{�����%�_��K�C������9"�=:�HZ#x�qIɵ]���ZW4&����@ ��������&��ܠ�s5a�&p����Mz�-���)���	}��/��D�<-oN�o���_��s�ď����������qӢ}S�S���@��.*>�B��C�ú�-ܧ-��]��}c�Y{�b 4�*#HN�ga��$m��nvq���q�[I�c�3����4�1m\L���d�A:�*g�B��}~/ke�k��G�<�/}u=�Yo�p�<�o��mq��زm��:S�f���j�m�m��m�6[B}Y �*��{���_*��ZT�ޟ59�l��U	�0Q�.
'�!@��s��$\��t<>����s�I�دǚΫ
+�P�Ӯ2=��֯#,���m����=�o��jv�~{X�]�V��q&�^bz�IJ�O�·�O�=���������r]M���;��=L��hd�@�;/��ɻ�
}�����R��=�>-MҞR��;��b�+vD��A��0T㢵��q\<�X;���1���ܲx��[�J@��W�o��*�t���P���%f�i�F�_�~ׄ� h+i �c O��6�^��6���H���I�5��Y��r�I�7h�5
������9k
�݈"��2������ k�B#�J�3æ����5ג��eܚ���o��1Z�	`�����9&}�L�����d���H#=�tZQ	[���M��zh��7����"3�SrL�^HP������@���)߻?�E�ƒ5�»W�m�
:�B�7\��^t4Hp�U:*�*n�4��K�pPv�ԅ�=�l�^�'�kρI���?�, ��f�,�ܦ���I��m(��D��.���j:Yf	��*̈�PYm؈t]x �Dh\�.��ń�S�܁��1C�� 2^�~��_1�Dr!��Na�0(~{��Ʊ�Q�[�;��{/*x~�\]	a���։�TL?������e�(�/J��6�m���׵{iu\oZ`y�D�Ee���%�B� ��~?�XPf�It�-]�}
�h�v88ο]e�w/�|Ў�eW��%DYRJ�|������Z莎��8T����ʭF�����DL�́�g�It����������n�"V}a�y7���Z��@��K�<n�kK�'�6�9D$��x��X�_�Vk���U�\�l4kW�5ںe6��YbVj��\
�E��,`p1#�,HAz���|@T�g%�a��W��E1Te��۪���2;{�r̀~8���y��1�>���.�_��l�gb(��	�$:8E�ZM�'&��7i�����<�NU��O�4�@3'c���k�F���U�'燞P5��{8�~I  pbߍaO�K����lu������1�g�������nj��������<l�;0g�3�]N�ɜ@�T��^W�\��xD����I4�i^C�������x��,��O��*�p��*Om�5�!0�Ǳ����r�Զ�A���i��/�l0T?�R��-~���o���d��HLi��Ҩ-3�d029��k8�0!���	p��7-|��/c�=�(�a�Y�s3��6B��>i>����'� �.g�b�>!XƋ�!������S�b�p�0�d����C�;ϥ֍���9�����-�s��dL�!|���L�b(�D�(@��7^��������&l5x h����W��&�^��p!ȗE�y'M���`I��~Րf5�>6e�P'7�ֽ]�}��;�Q(���|��_ +m/M��ic������<;�\����+�cF��!�Ư�R�Wcżry��LeP���3�2�Q�>���[��+�F,5� {�zn\���sx��<�ya��t�P7��V����#@���EY��H�T�s���;���K��cNCB�I�R��y(��<<7jQ3�jxP���yh���tu����K��϶���	����+������/V�P3��}B��mP"��S���cu��]}�^|�u����n��O$��<ZU\�v^g���
��D��� �}s��3J�{�������顩��B��}0�1��.��!�;a�ɺ=�r ]�Ko�۰P���� ��]�����oWF,ܳ����X9'�?�e[l�����X���y�Њ	��G{>�WOwť�:���ŠZ�z2�d3ﲖ�,4�)�l���7[PO�a���便L��,{d���iis��tm�h�0�P#: �'��.k6,�͝�YH	�k.М��[�����_^x��*�\bLt>/�Θ ҨɮQ��>R���oz>��z��0Z��׻�`
B!��5~�F�z[Δ,����դ}`�����K�I�8,Vr}۪���h��B�]�<���^޼�{1�:��/.��×7����t��t�UnWp�r�mU�F���a��5gC�sER�+IZ+{dd	����M]�k�������-*�,�|���UID.�&��62c&��ҽ�e�+�_lr#�Un �k(/cs�!�8��>V6��۸�x�I�J!H���~��l�l&� �I�	[ح�ɲ�S�B�IM�+<��mAN�l�n���3�����H��J5r�|x-�����`�h���D��D��)j3o
����1H���w�9��Q�D��Z���B ��,�Oz�#,y�I��Dy��,9b��	}���z�����W��.Dn���n�()5D;{�P F$?�p�dZ:��E��Q��:�1��+�/�bk������D��}�x�����A�dn-�uC1�m{`����?�)t���1V��3˹	)IC���tB��*-p�s���!Q	G/��,���E�;�^7c�A�C��� zQ������lC A^"8���)y��Q��0��/]��d�Hu�f(1�=q+U�*��S�.��ڴk�}k{p�w3���ue2�(�8��_:������S��8r���<�&�"��1��l���t֭)�I�ʢ&��*��{���o�?�.|� ��AU$#��.(=g^��;�����;3�Z�D��I.}3|cLbrx�����e��O�չ�����n��ڦV�k	v�%2�:|�!NZ�ӠF�H���'�N�+�q�4QG���+��1�Sh��i��"�`Ip	��f}�3���G����~�P�� ���aA����mx���k�~O���=���8|:��� ���[�R�t.p)kj4�n* �z�����tk���h��0w�����u�\�G�=)k�ySa�x[�Q���
�V�ڗ=d���#`q+�ɡO��k�:�����3����$�jii���=��A��A�:{�m"G�½��=B�Hq@�غ:z�1��l]xW�����ِ����p8Z�
�jP�)OّC=�P�3_�&�&�n�I5T��Q���x�GL�Ƒr/�JL�<��=5�,�Z�B�PdN�|�(K��ʍ��y[���c��H�	�_u���_��Z���m�(�r�Mn��e�GF��#ѐ��(sN��E���m��G��HR�i�*�������h�����I^���-�U�W��&行ǊO��-䝟MrE���m?��'MN|e�m�N�N&���?F�
m�Q���r�pi>�q�����Zϡ]���0�0��=EO��p��{�N+r��Y&����	�t�M��3Qnُg����br��sX�ƗhA�ׂ��3�$?���KS�մd�m�%[��{��jm(����j!�"�;����ʏ����+\R�Y��re��DV��?<���mN�)��ut����߰K��%�m��$R�䩍-��U1�	m)�P~��Ry��7���5T!Xc�}� Q{��lG��U�G��= �U��n��K�!�%��,x\�BA-�K��� �A�j�笯��r�I�ˬ����l"|֤h�a�]h�J^5�S�ߪ<��_���[x+�K+y�,���ؗ��y���C2Ǯ�Xy��k.� xM�ꌭ`����@j\G���x�g^���1�E��"�ldu���nƇ�����6@)�׺�lW����^r�H�F-�;C��刭!6�49m.�I���<j�4�9$�O5U��V���������d|}Jإ��M�����1���w&>���Rպ%n�x��j�ѵ;]��H�#f��)���(M�f���@ qN�_2���u#�@�TF���+���㫼_�
�7���+K�ݱ	ǭ��O��L�&����&OSq�d�q^�؆�E�]�������sV-_p_��x��`t�G���jE
۟VEִ��I������T�4����g If��A�h���|z�C�-��^@���z&q�`� ������ـ;BӉl�V\9�Ƽ�`c�0��=6�	=e��U<qoG�>�Μ;�1WM�$gIO\z��U[��9�A��324ע	o9�ɠ�q��e���t��Z�k���Xڍ����#�n�5z-]�C�
6�`�s�����l������T�<�SvH�5weaP}CjOp�����ųC���93���-aOy�YQ�
�����	1�{����o�q�re�cPƛ5+����A��gR�ݘ*��(��F�`�	"/j* _� ��v>qr�}"C����.c*�
u'�`�3�v����,�:$�X�B��ү���덳1Jq-詊tr���D�Zf�EJ��+c"�n̹�A6���\��}�`�Ҿ9�̎��)I]���O�X���)'��z��K���f�yE:#� ���z��E��uLK�x�KC��`Rg:P�,�N�y{!�u�B*_�(���P�Sg�⊷#Ŝ;(k��\4�n::7S����Z��>�$-�[�����*�E�;� �sU�l2'~ߏ�;�Y�x�0�,�����¿��Xus��jZ���ڴ�X�S��($�y��E�:(���{K��b�>�V��Y')uU&_�@����K<�� ��ZЙ���2N����:�2'8LO����"4��@�?�V����N��?:U8�t���8iߠJ`�[$E��J;�&��q�K��Y��)�O�\2y'ާ�֮}�����]^:T���cf+6��E+ò�,��pT��-@���t;nE�ςu�����H���z�a����"k���ܜ+s�*���I̮���Y͉�\C�����}	�D-@D5�($�
���ɗ[Ql�๻��^�=}9�5[���x�+	гl��,��3DN�0��/���aF@�i��)T\B�Q�g�}	�d�X��'�!������ÿ#�L�|+���T0!�x�t��z�o�k�.�E�<�`*?�y�^��b�-�+,�1�Y�	{)��F��K��˘�U81�|^�"U�M��K�5'�O�	�Ҭ�����˅.�zey�=�.�I�\M��d�r�A�����Lj�	���;������7ݡ��b�������I+��⢺�"Fr�"���q�菒,'�Sj]���P��Ԫ��#徧)xl�lo�\�(�C����jj�^�?���Ƶ���i{��d=ܾ��jeo�����p���O�Hy9�Z��)r3��)s���Ph'Wr��?����4;@�����U5u�}���5<΋6@E�%��tʭ��Ռq��}�vǁ��%H��CA�+*��CG�a�q��
*|��.$vI�>~	�����K-����ׯ\�l�-R�u�h�֑�D`ܾۉ�0�#�ȝ-��?q?z�"��=5
�Q�<�~$�H�j�0�4���`�B��V<��̮9�mdE�М�,�"��&�Mw|!���4�%�V
)f��N���S�ն��}�5���>�Mbl���K�N�{���&��|����k1D�@6G�K�����q^л|*o�]e��Be�IM������n�n�YI�F\\������3B�*`;�ࡤܯP���ƣ)�s �0��z��H�}!�Ͷ�<:���(؝��ٹ9\�(v����c�2� �7]����8kx����磀�����7��r��)��rfe\<c�ԹUMI:�a�Å�|w,[s>/^�'���1�h��+���o����}�A��l��2���;d�iع�k�5��C1B֭dxp��r�a'�I����/��8MX�ӗ�i0:Pp�r#|�9x������m��o�29�5ʆB��^]�~|�RD��iQ��+k�	�8�d}�?²��zwŵ�,�-%)<i���4��8��}Xҩ�0U��ѿ���˫b�FwVak�K K`?��s=
���[�qԔ�Y�sk��)䄽�R���!B)��2�'T�n��i�判a�g�vF]��wէ�/*z2�Hd���t�Qg�������H�nX4/��C�@+QMeL��ԗ�<`���F*���W���-qJ����9��"�ݑʔ�[JI�CY��E@�H¸��m��E�~�U��I�1ht>�ۦ�|�<1~k(���rM��o_��֋�� %`HP[��yuK��ǅA�*9B}�����vT����؛���г��n �Y�\R[�rO>����t\a�ā��V���tW�42��1�e5a։Z_�X
�I�U�Ȭ�be��8��t�Dc,H{
�΂WX����������I>�$m��F�دo�>��V�r�_4�R�-���v%��G�y����il2���F�=�Fg�t2	?���{M��+[��.F	LF�\Q�-�����C�<c�w�*������?/+�0�7�hNa��Q�����ͧ�����з�̠" �����/�Q�S~v�fE�	Y?C&f]���2"-��#�g��{E�U�@��CU`����WT�����:�:��w}�	2��	��s�Wx1w����>�6^M5$#�1[�k��j�������C���$�sJ�:)B"�Y�a������Ywb�fA��I�m�-��}�e�ɟ��8Ƥ�k�n��@�4�����mb˾&�=T#7;s�yԨ�����7�m(�JO�l� �
���B���Ϫv|��m ���Ӡ�,lt�e�`S���w�_#	�Ue�����r���gL�2�Sk��-Q]e���8pn*(����2����bc5:�ɮ�F(���@��ts��ݕ2et��@L�5�!��(a@�����j�z	ZrFH$��F=�-�i�i$y|4�=ڟ[�3\���	�,X�R�m��&�%��s�:�Z�g��b+.��ɖ����w��K�� 7C�n��pe�	Xj_��Fo=�����[
�$:u�	x��qJ�Z�5�����<q�GӘW	]g"�09�-�����T6���W-�i� yR�Yi�|ky% L,��^Ӥ�*5�� �6���ZZ��9S����v>j��KԵ����%��b������[�>E�!�Ĭ&���~OJ���YĿ�74���m���_��^*���D�X�Fa,>���{�5�U ;E+@[+s�Rؓ����B�o�vW�x�k	�KdK�_%O��d]�+�1�)����9�L�I>F�e4��ʪ�L�n��62ina���&@�6K��{O�I��n�3f�}?��0<�7��h�)>ğL��z>T��UM5�/��"�|�:���iW*��(��#��L�[w�a�0O�5��b��⋮�tU+"�)��S�S����|�|��>Gn�AKX��� ��1�E�J١?4M�V?� ����2ߖ�F5�Q`�����=��?���bo()�	!	1]�3��1��D���f)4ULW�)����P�/ڂ[D+��*}^韣L�1%��go��q��^�r*�R���x��<�妶V{��.X�S^�v&����Kik�����΅�-b��dx#�L�&����c���]��������M?�2 n*]+ف��L�f��ₔG���������� ���!c;�a�\�s��/�������O��LL<:8�l�W�p�dQi��;r'��(6u^Q�W$��W8Q $?[��8^F���d�$�R�`X���s��+�0�b8ac����BB}�R���9+|(T�,�����:��?�w�l���S^�q�4��ؗ�`+}��h*niс���=j�9z�L�F�OH
C��ʽ�Ca��Iu?�������N��ů�_q^�4;6�H>t�^^~2�ɰ�ٝb��ώ�DG�Qb&k{��IެV����i�5��a�D��h2���v.?gl�-�J���]�=w�TŴG��h{����{��cC�g�\y\tf������<�Y�p���L��mQ�LÓ>�f��|�����ƐNz�ok�3#���7b�')�ւ��*Gj�x��"��qHb�I���o���ě���H�f�I��릙Y{y\��20`h>��}�i��6\!�TS��!Q�K���5W.��T��Ϻ#�EAmw� ��X���K��z�Oއ?NT	���Ӯ�'�m&��ή�{�8I�Ծ�;?I�=lT{6���۫����V���圆B�l�r�Y�n
���������A�f.K��� H�]�vFO�k�u��$Ѵ����+r�
$Z+~-��yE���Y$��=��n��H5�[�T�9�,������
�>;y���M����Jx�dO�1.P�L��5ы����9�t��<�ݫ	��z����]S~�Y���}�ǡ��|_̈́!�U	:%���ʚ<y���=��=Y�O���*3�����k�n�n���rm��6�J�����8��~7r[�9;�"�@��W���4T�X��%�? &�yݸgD͙Ơ���\G��%��Pa�3|B�+ۑ���c^���0�r�s,nc?���ff+5��i�U��9����M��p�"�M�s�e�"8V���7���3%�T]�v�e[�'T�As�a0ډ�����-sl�����"�����I�	s{��^�'�����T�~�aD�������v����pwÄ҃�DFi�Y�C�mhM>�t�<���!���������ӡ�S�I�m�]�ȾGb�	_t ɜ�����Q�J�Y�%"⃺�����w	�����͉�b �r�;w	��u��5��+3�d�)/�I�rxĂ���P�X#�`��ǝ|TL�x�'u(�ܔ��B.���A0���.B୰�S�WP0�eA1�iI���"P-�.{��Rw�B��i]^">�M���-{�xA����c�dM��L ɉ&�ıl�z&gK�zTb��9d��E�ڙ�@�5E'��#2*t��&�����]EܦC=�)}F��AEbP��	&����4b#Y���e`��BZ�ʹ����Xv o�^IF��'=�^�B��R�H������-l���������D-F	���t���]���3���A2[��g������Wn l�~=��N���nS)㵧��tr�&�����x������tT[�ݻc�=*%�{|g�!�Ȅ�����&A<�C<�)�d�6�oۮ���2��>D�Y��|R�;#�v�~Iu��/K�Es�K���8�BC��F��¬qJ�ͯ��
1�cQ~�)�VoE��o��?�$�죾Yq� �퉇y���QV�;Ã�]������L�<��~�R�U���T~T�m�h��:�_�d쇰J�O�ݼ[��励�;��{s_zL#��8Y���^�H�[W5���{$�/r7��xH� N9a�Om$w�-*3 �r����20y�r�C��!~�e!�9�����h���֊.RZ�Z�r<B�Rj���̫/�?v�ɐ�ה���hom�v)6j܆�7��,Gv D��<,�_[Cv"�^9	K�PEf���e�I��'T�5Nv���{�@�u��+e�lP���
�9M%h���r���"��^�l��{/���-J4Cm������=��J��٬����~��^Z[���9�^��y�`���D����T�v�zJ�5v�|�]3�m�����ӭ�q0�>㫠�H�fO~�b=N� ���΅D�O��^)wr�[HV~5�f��p�$�XWB����>�+�)�1"��5Yp��r^���4�M(md�`UmE��}�W3/Lh�;D����E�@����/�Y���k�ͅ�1y+�W U��^>LD;�΂h9=��	�VȲ�A��2n���0
qO��Ya���.\癫��qߪ㜋�&�Þ%ʾ,�X41:��/�+��KlR�G�+��)�U,��,*/��� ��TX�3�pUe�d'Ab&5�J!�/��n�!EcK���01w�s���"�����k��ˤ(�e7% ێ�Np�'\ɤ� M[]<���\�iߪ���A~��12��a	��������T��\%�[<�}@���UI7���E�?=�B�����qa�^*Fܼ����Qݜ޳�>V�^j���9�8�n߾e��#Ö
���&%+��-P�;�D���C[~+�h���B,����i�b ��^\�^�}w9�⯞2P���0�w�6U������7v�E�Zyᗛ�w.����Lw@c�+�/Ǘ?{�>�P˦����΄:A|:l�[>y<_G�	I�e�v���wzK��?ߓ��Dg�2su^C�pr�Nvj�7/�+{�*]d�.� %�;n�Q�'�Pp��Q�gQK�7��wyQ�Mb�:�QË�=B�>O��(RNΣ�mS�5�޹,H}�]b����bT�+^j5����ïT� -�8�j�UMs�t��><��)"�`Н��;��	�v�?"f2|�|�"�#�c��煞�k3�?���5JC�Z��F�;�2:���$J.��8��Ϫ��Q��=|JСm0PK5B�K5�.Md¸Q�r=�dNo��M�B�u=�ݮr@�T��%k|L]�us~�7)�3��d�+-��#Y��H�7nA������}�[�����j̉�@�(��n�~���
�3�>̪Do
��|	=^UʝP��Z0�]�w�
�:z���f'��l���K�&Ǖɾ�H�=�+��m�v9ƞ���;T|������)<�} �j#}OU���1�k�+�U�����nS�c2>�k�lh�G�J��-�I�1�(��@\xY��b�`�L�����᳁z���k�pU��*SE;�}���͠���>�g@SϠ�+0y|�����io�?������}nu�yN�ӵ�;�ށ u_߿�#��3��<, ZJdg��[���GU~��Z����(���at�d%��gZ����bn�8<���QOMT;��ҥ�x#�C����f<k�&��B����������F�����.K8�.|��|ʎ;f����
��3��.��F�?Yׯ�D��[	h���s�&ܷ��K��֮�������
�590�Wo�_�'ꎞۭw�KQ�R�]&�����/"]�P�j#<_��{����8�w|��}Vv��� ̈́V�u���'��GHw�P�V`���^5�'N�xG�-^�M���!7M�Ks�0��΁��#�c�����} <���#�c+����oR�i�yK��&/J
���-eD^GiT��;XM;y��W��|��о̖7{���`{{�)�F�$d;|�����I� �l4á���+�YR�P�aݔ/��/(����H��}�9NT�f�o�����e��7]��Ƀp�����W�_.���>�A7��-�$�8�N}�����V�:Q��Q`^݋uX��UO�Of\5.ǁ<0C}���gf� �>7DI�0T<%���8�Ķ(�L��BG�D;�&Q����-܂��R֑&v�
������ �䊲ُL]S�Z�i 
����Q��������I4f��Ŀ�����ȑ-;����	��ߊfe�Qc��~�$�� ��o�^F�?7�S_1[5�}5�79�FC2��QU���q<HY�'r� L��,�����ϖ`�����u*�{9�$��AG1W�Κ�rA����>��b��L��5!N�+�X��{f�ԕ �%i��8��ٲR4+e�L���(�mpNm���i/︲,�1?�@�>�+��hP͐I~e��cXcvV�B\jC���rE�/�5V�1X
��X�z�����9Ѥ�� =�78L?�2>��w?���g�D}e90�3�\|�w�D��_��O�����Vh�t4s�~ۅ[}���pǠ��V���7���9ݖ¥f���*-�Q_g�M�Ш_:�9�+�ky!��l��y�e�������Aneuw�8&%[gz���'o����fS'�I�G�Z+Ĵ��ͷ\Os�����h�� O�Xg�I�1��A7*
V9�5����Z��x���1)�8y*q��,P-�J���5�kV�؞4�z�Mq�gu�V��Qj"O�R����J#K��*ￛU{4�Y!;%�ƭ��z�7�D����|!�N�[�Z{���y�1j����x�9�ђ0�	;��Jp���H�:�f��OI��Ǔ	!���n_�=�#n��89��o��"�0�#��E#1�ൣt��)�[�	bw�����~�f'�,����� G��e�%�(��G��	j��Ȕ�-��j��L�����c����ػ��3`ʆ�"攠��	��2EI��q��`K�@!u�� ���F�5��UF��6U��6G�\ZP��-�W?����%�wo
�S�&T���I��xƠ����3;���e�U!�<j�ƨ��	��}:)��Je�.�l��.ҷ�F�R�M�X;#1�����Oe����U=�0�B��3Z=��gQ�y}GO��s����������'Ӂ���A}�=�����7���vg����h�
��zM_&Y=ލ���?6�p��;?�����|��R�pE���P|L�pYB'O������k�פ-���Վ��b�C*|���F�]�J����s��������1�����\��C�⚤8�'<�)栦}���ihmX�u��B�����@����gF�$zG!��UW��!�X�Œ�ӻ�7��In:�¤h�\�Ȼ��"��d����O��`��K�xzB3yM�����Uz����E�sW?ɪB�nr�X#�W挘8���۠�3�x�xc[6kJ�2�[*�DX���bl�.�O�=Θ�C��D�FT�I[�^ۄb6��e�I�/�C�߲A�"��F�pRiX��L�'�躶Oc����8ߌ�R�R.#U�s/�mg>���A��3F�]��qԟ�ӱ�/��;X$v2��S%VO,<� X�K>硍���=�:����L��K�"> �r��J/Z���X��/̐.�-��iܚ~�BC��hfC�3�9��z,^�MT2|A:�����{�#��b�qV��{��1���[�8��m�'f�������c+&���9�^�!��-��~�ƿ�Zӝ�_H^���`t��}fh6��Z�\G��z�C��D�������O���r�ڪ�I�n����U{����.PU�)]�M��{�[V���_�?���8�"�s���DQ��{���S>a��k���<W[�����(�D9b����nsk؁̓/����:�hħ����G4 .8b�����db@c�2��A<mu�1����O�,͗�ɹ B��e����Y��i?uY� ���+7�s�?F�#��"��gȳ��Q�K��Fl$�fBU�b'd��4zq�s]����	2n
�A�6(�ЅJf�:*g�zz��&���GF7���ȈOd�j���{Q0~�z�?ӻ�zOD��p��F˘K!u�վ��v�T�OW���8J�lE@+��`�2�z�9x'b'67v�l�� (�,����̃E�������`8�����G:�1�o�4���+�z?
 �q�d!C>�K>c�%8��.U�6я��ƂȀu�a��맡w	Am�-%���R�
�k&I���4���9 բ�$
hn�E}�g@�-V�d)�Q�d?g%�bT2C3�D�h�ہ-�Q^L�M(d�*J8�Z��𼬛�u�as��Rf>g!�v���U�夲d�-%
[(6��(�Ao|�{����F��^���g���Ln8P/}s<�^}�$h����YJ���3�Ut�r��m���_T���a)Gwf�t��M�h�����{~�v��z�p��cڏ{�U$x�_t����U�&��ǩ�]<4sPjZ�mr:�Ť\&S7��K��I�������<�S�~u��<;���3v#2E�##���bV�cGѮ���-��(y�6�i ;����41'͑l	��3x3�@�������<J@5�
�l�,�'�����R�)�Q��]!�/Y;x?ߘ.��xW��9F�N:�i�\�����YD��]ӗ�"ￍ>���=� �ƒ�� *6�<�I��9�C<�#D���/�/�o樠-C�4)��Bא��(���|��5**Q!u�)�B�H���ռ�L�Zj��������gv�k�j��Ua�[:@3���%̝���%"���yB�����ڨp8c�ߝ�}GH⹂��k�v���b����fJCs�=�!K;�z��&�xӸs6<y�m�p��G�� �����w�n�Wǟ®��ՠ�u�s)��E���̗����z�~j|�9nB0fMU�Ev�	R��3��������Ɏ�IG:z�*8�,/���ՙ��,�H���k�;o�|�����;���C��+QV�M�f�ȟ���%c�QԺ5�����'p�m����)4��{�Y��d�ؙN#�����.x	ҍ%J(���G5_{P�@�u��TM��fZ��θ��@i����6�6B�(/���
l��K�$�2$pn%�������1�?_�~��J�D�����w��.@r
P�b£�]�ܲe�+Ol}��w�ւ�0[]#WE��O���� *�՛�L��0�M[jS�q)�t����8p��TZ�r����
�T�3�^N�葠���V�#�ӆ�m湪��0�'!�:{�w~Dmd��ڎ5c�?����O�5�ހ 3j�Erw��5�������O��n����x%�\t^�Q��?!!{� T$�EBVO�y��M($m�Cb/��o�N��W�I��s-X*-�Urˬ��xu�O-�$z�]+�]F��>Hj�8W�r��0;�S� 6U��u=����_R8���N-�/�������&���Е�b�� ���ۢ{�к�l����Df�7�,J�g}��Jr���� U��!@� �Å��e�ߔ��<�\g�!�0T�4C.���6�Lw$JI�i�Z������ڱ<�(�)#�Y^������m��6d����X�/L���I����
�A��1�5~���}�0�YY`pˮ��[a)O��w@:�����:t��\���.�ƫ�ˢ����24	�
,�*�]��X� �v�+C�+W�(���N_bU�b�D,|�\�
��1p����w_����̘)Vʘ�v]�9���ߏ[�����=�)a��Τ��M�f����!C���WL�v]���٤�� 77��2,N+,�Xvh�*b��!G �	���&n<�.�
>X=ޯ��ji��:zl���x�;�m�#w�?�~[h'c�	��k��_�Glܳ�bLz&��ŝCE︻�%����Rh�Y�>�_�LyK���u�ҁ`��4���m~��:������'D�{��Ul�ănh{}�5�e�D�$-*^8��n��Q�iNi�D�\p�\�>w��_�~�^��m)���B{˔Q��3��H�% Pf0��O�Àa��h"��J:VV���9������X/g�sY�K��I%Ա�>���Uq�VO��0�e=�~םs�F
���D5 tw�u�Hd�VS�$M�ړu�
NQ~�=����2���d���~�&T0�+�B<!��=�"���H��(F?Eu�_d~z@梮O����'q	Y��^m|S�I����)�qD"��(�h� �E��,�����cx�qN�i��L�{�Y�~��䳀�ÐG<E��r��T���BZ
9��q>h�>��xL����7X���������Ջ�3/�3z�5�X �4�k�<���O�H�ya����ɾW���������lDj8�$1~V��B���D�������a)��v�Y�;%�_Ѡ�X}i�7��:��#�}�3?�����%Y?��C@v���V��0�m�*��
n��S�6�e|j����Y��Wy�����-h����䬥G�tᵝp[?-�^�Ei�d�ѯ��;�Hd��>!�0#^Ӆ�Ii�@C}�^� g�ʚ$.�ι��K���#������ę�Pb�}c����E�<���H�	1�#c��etޤ)~Dnf�FgӘ�BN��!E钭�l����g����TT��Uq��e`��+�n�>ΩJ��'P�g�e��v��Edi%3�O&Mi�Hޣǚ��X�r��:���l+�Fl�WV��?�Mľ�AaS�Iq���݅�
���6�(*�l�YV�E��I��q��ײ����	�H��VN��5j�ؙ"I㏣�Q��B����X�O7X#�i����~���w#j|1g�:��j`?%x��b��'�r�	���b33�X��G�p�81o�ϓ/+,��H�#ΛO 4�t1~������f_x�Z#/�����d�S9��S)4�R��C���DqW��ٰ2ӒߤM�Qī\�L���-x�c��n������ѕV؇��\�L0���� � F#+9��\mKyh	/�� �^����{0q��4D+*��q ���2�K1�k^�����L�7�qcž�c6��n���m����D��5mA�����>�3�{*xB`.P�tB����Z���|�]�c�t.�>�Kp?O��R�l+w��v��-��b��ȏ�L�ƚ�X���R�r�J��\/���v�>L2�}�8v�&��^q�Op���eha$'�̊k��\�]� LIo�_+nW����������ʸo�y���޳���B\� �)���{��`�V�R��f_�b	�i�'��g�����@���u�lH�h<9{��k�%�����TY'=��Ao�'<�B|M�4Y�d�Y�i���7&-a���n(��*%ۺ3����5~Tgh�g�b�K����&ܵu�X�w�}T���)K���(P��0
V�_�Rx��ȴ���l�Uy�)��Gn��3�!!b�Lz����,j�P��MB}]��b�<�;��%�$}��`˖��prF�jx_ΐ2U��vPG=R��(�%4���ϞD�}�,Ʃr�/cM���;���$h|6�f+t�S��q�{�'Gv�R�YQ��
*�&�Z��
�A!;A������;�.3�Q���P��,����v��|�9hr���m��!#�5E�
�?06�p%��|���%��T��2���OG{�'�l|���y�Dd[9�bm�H�ؚ2K'�1�~�Q�e��Q�߾c>��I�Da�:-i��$ A�,A�M�`G��]f��E�RRd��<�l}{P5��$)S�VE�����/����\�Ǎ�aM��^LJP�����[�ڗn�oΆ����x�) �GfFM�F;-�0���'e�z�7J��j �^%	�T�9ƸE�W�r�.xtZY'�����ڒ^�hmH��Y⟟�{���m0��f��ġ6����B���Zf*)��DjV4ow�k��և���4�>f�b��P63��9��~��~J��ˤ�p�a�w�"�c"f�|�E3W�e�?��ױQ����q�vɫz~���{����*�3�^5�mo�,3�w�=,���rN���fo T64x,�N��Dm�G�/�������F��@u����Ѱ�?<0~K)�!���ׁ�7���tӧ���sc3��H����h٭����7��Џ44���u�M��'�%~\�8���5��+t}E�v��a1��AF�:,�0 ��A�����QD�gRc��%�N[��Wޕ`�*�a�&��Ё���)H�G��C(2E��jo\2M|m׎z:�`I��s�1�Z8�24�Y������Dx�XhO��֗���r�S��"����z���t��P�d���i`:��b�~�;f��(��yvxM4f�SD�sr�ʁ�������	�D�c��Z�XS�K�Rë�}��2�Z])��x�a�O��O���Q�3��̶\x�W$������Lѡ��	pP���A���v��HN��]x�*�6�����D�b���Rd B�+�.�k&y��3�ȷTLEÊA�(�D&����Խ��%]O��21�JV�'Fv�R  �u?iq���a��?�$m�/Er{���<��p�(}�{�Lݗ��`B��2~�$���J�j�DL�U��iA�O{5���q�v�qVP���~� �ď����>ao�~�{C~]��8���!=m�����)W*������������<,�i Ѽ%�[�*��ID|9C�Az#���p����*ڹԣc |xc<:��>�a2|!�(J�Dm��/	�m��^��F�%K� p�d�������n��g1���vc6-d�_��t�%�����f�S�Ԃej�R��q�[L�2�<��9�8~�Qˎu��:���R��<��o�h��%������CE0%X�p���� -G%���9��#�^V��+LOΊ�;�יp�]#���{�"�IX��a�H�M��9��p���\�/]w$�B�\W�E�hʌ́�PpM�5~Y5}%Cl��;9�����?�A�-����`SC�hJlM[�^@q*�D�#)sww���[n�)�M��,
�1}<�v6H�2���f�g�Cto��c�b�lY�TS�x�ǯ͢Ϝ���,���İy0_�I*s=�� ��=b�)����j�[ Ew�o�_�3<$B��@;��
~�r'�+Κ�Q��m6J�����OX8zN�\G��"p-4Y����z�se��i�����8VQ=��;a'�<��"HY[4/X�a�r����1��Z�"98�������糉��F֡�z4�CQ4��$a��$�C�R�o���9��è��S�$q��o9��t�^CU�ӆ�6�;Fw'��#�x~4{����Q�̢���@���9���欥/d�1��>(��]7Y[�Ek:c^��m�L�M�^��S2ǥ�?���wDc�nOL���޲�R��Xt��ȶ�Ì�ԇÊ�։���Z�}��$�?[�.{*��aB�c84�ނU㠞8��{3�J��H�u��&ʛ����"��=ʸ�^T�ed%�w1i�j^�=��3�x����[n�Z-.��,�����Y�������nٶB��\yq�[m�vq���;(Y4�;���A��q7l��Ĳ��O_��T���R`��0N�=1��k0���R�.�BN���|��0��6c,�TDE�؉_��*���T� F2��T(c��g���-5�d��\�y%z)���&+oA�4��Q��N��U������7�t�k>�_`'�	U�Bl��Z:q }�;1�KWM��������Z��Q&7��0�U8;���:J�)�|�^� �.���
���9<2�E�2��\�W��V��V\5_���AM�E[]	+S"V�ƭ�O{�m�ă#E��� �U�0� }�1�W�?���`��R�.kwF��j)/�?�#-kgV*��F����bMO��`���}��ِ�:7ڦU=�;��&�li`À�nʠ,jZ��&���jK�E�uY:w�飫�{r lbA�V��8f�r^;�,���L/�E������=��vS��S��5.�� �{7�)�Ǚwܥ:@�a�ҟ	���H�Y�r7?D%����UdגOb��B���Ô����Jb�uZ;����8_f=�As�ͬ��'LZ�4��ۙ��f��X��XG��_/֞�Êؕ�%��$//3V	
��>t�R���������=j�O��P�t�"C� >��y��`@�v�P�Q 3��Yt��w�x�T�J�p��t�&��~s����}d����ƫ`��ױ%j�z::ɓ'f&pT���6I�(�rr����T�;������� X��@Q����2l�H� �ֹ���#'�Ր���(�������t�_8~�R3|�h�99�``'�|uOP'����M�q��z�AC�cZ�b�ɰ��.�^������
 �&�o�}����c��̓S�#gʺ��I���\�$�q*Jx":_�VLGF�z�0��H@��-ske�pn�����/ႝ+.#�/(=����F����D���S�uP�¬7��Bc3t�hVz}�|sa?������m�i�������l��"S0#�kJ+�b$G�e}3�ƻ]��o:Z��Bj���k%�/�6D�	�M;�V΢�IQc��ڸ��q���`��)�o�U�4P9���FH
���E��r
K��&��Y�%�5T�z�%����ã��e�Z��S��I�4���9u��!P ���0���*��m��~�5ʽ�S�z�B�mk�
�Jp���h�pG��6�u�<�Q��*#���M?0 W����UGD]����b*��|�1r C)K�m�������wG?��U2о���,��#Xd��FT��]���bGP��Vg��y�I�V[��(�4T�'�ۧcPы�j��s�Xrc'�,}=�=��c��&5C�~g��m���<�ש�c`�'!@��ni�l��vۍ��7��<���Z����R��S�ه�f������ ��vH\�~l�OIv�꫶�� �6"�j�"�Ҩ�r!`��]�<5�����<�lBk��`�#&��\���B 㰸S�S�P"���^��{� M�r���b+ǂ�,�`��'�I�{��	`;���t��D�YUѭ'�7���|���~=��\�|��ݨ�c�#嫚�ͤ[�n�Bz��Oa����d`�C� _������з���0�%R~L�\yֹZ���O~�����sk��vK:,)ܵ�QC ��G�$�u�yv�X���Z}��b����36��d ����0�%N�ƙ���qjAcvu�6U�%���[��	N��ts�r��Ok����oK�Y��@�oF�\̂�s����	'^"�/�5�N��9c���z�A?�	�oW��{�I��g��;���x��E�1�Z1��3V�L@�O"�-7�(S-��G��Cd��G(L�4B����x1�ָ�X?�g�}����t�O@RXB��W�Z]��V0��������a0�:s�U1^�N�m�`�.��=�;�dM<���ż\9ѥ]ktO�!�8%_��zP��23f���?��R�0����U#��ӳM`,�~j�~T���
;��*(�/��������ٗfR�/���y�%���4�#Q�>���!�����[�:Fgi$ڂ.n֓ �|FkL*N��E"��۸>�z�J�3K�!�F0X�U��"Ԋ"�t`+*�Jʾҭ����IBzµ��-�'�Q��3r#y�^*�@����9_8i�$�P]�0f�����+黣��fs��_��*U_��і��C�2����U��� 2�D3�H<0�qF���+�>�'Ʒ��H|�D/�&g���k�c�3��)��.v�`ڔbz���|0Q�3ې�� h=��'g����b�1 �lA=Y��h^v�Z��N��
��1��o����ߖ�w�HR�����X�=�6e����u�[n}W���dQ�����>I��P	�I����5��[={ZI����$4|�/	+��֨:`�X�����r�K~d�⡩�pT�ݳ������;�\}�m8=�>�H4S��R
%V�0�Ջ���W04sG�_�\���
y��C�0k�PP��f���f�F����cw�Ueu�?�&'/'��l.9�Ҫ ����1Q��0֠0+T�ז���_k7h��\R���Jn�x�оXn�8C�h�~2<8"Y��N��y��l�x�ei�Uj#>U�M�§�,^�T>a�e�NJFE�u����A1�x�������<}̾&��x�Q�Y���{;���N�<���ʷӸw��~�=S��U6	��Yo�,�U����< 2n��
�q���z����Ofh�YQ����ˮVz�^5�a�A q�5搡�}���˓��V��-����Qk�B����
�]��KOy�d#�B�{K/	C,]d���+'g��`��A���yԀ)�&ؖJ qnm��$r@�8^}�S\k�Q0�-���Χ ?gQ�M!�ƿ�R�K{eU�9~��L��׹��t�Ʋj��*JV0�I��p�N��������E��$�����o&�����e�����[��B?W]
�xfp@���|ֆ^���ԏ�Q"/em��
��ѕhI>$�8�]�X�)z�N�zB�����2�Z�����j7�����m̑׸�~b$"�~��J�wC�b����͂�6���������41�H�2r�k*�r�P����Άos�m4ۖ0(�OZ��rD��
�tD/zx׺�ڥ�R�R+�t�_�&y�z�©4n��$���ɮ��ChJv���I�Ρ.<��q��
5�'�K4�� ke5�4���???��:z�)˅Qw���{o{V[4ޠV�i���@�P�s�̰퀱5ʂZ�E����A�A�c��/4�m$vt��p2s�q��^�>��S�<��M.yP|s�^�������uuS(�ȵ�6���>*q�c��eu�Q�A���62����unA,l�EK�s�.�։��+Ѯ�1�?.j�b|H|�BcU��=��6�R�����L��V?p�I9OȊD�OenŜ��N�N��ND��Nf�k@"8��E�k�{�j����D��^1Z���c�m��AG������*�D8��s�`6	��K	�X�����L<T����n�q����bD(䗡�xr6혻N�L��LII�>h��7Ġ��V�%'���Ů=ϼ�	�7b�8T��[sV&k��L�;����mQ�m9 ��V��6�"%��f��al6��4A��Ē�8�w�',ƹ�q]�K��!k���Y�:���C�FJ����#G?����!8^]��Վ�X{1\�ؾ�U�b��[��Px�	�s^�����4�&�w�sTEK
^?�������#y��r��:�����Y���Q`�#��1kD���]���z�t[�oC	Yұ~� W��:��ΐ�͊A/��U�}@���e\T+A��S�Ed�}�x���m�Wlc'=Z ͅwùR�-����G�w ���̻���q�m$��l&��=����	�j�:�w�`�24)om	I�PHBp,[dK��O����i
OO/��wu��<]ܞ52@�$~�hU����/�H��Y��#×4�ȗ��w�ݫ����)���c=����:�ϾRtI@΄��GrG�N:�/�&ۅ!���+��:<�J��|F�B�:"Y��s���:v�>@p�"��Ǖƽ��K��������&t�z(�~��e�B��su�>�����;��=M8��-���zhc4�t�r��A��xE����~���\��/�]��>.]���Q.�<�V߂;-%֢�!�p����Ê��9�K514�enS��G�T ���a�m�]���6����JF�U!k�.���)A�Yp�Fr�=>7�&��+��jI��i~1I�!bVB-�R�m-��A���b��3���\���
��>�<s%�Q�؆à`���NQ0�lS0��a��>��@&�/�|Z������#l���#�:��~��2�5j��{�=�'a�9�[�ʻ�m��Q!kV��ؤ�%`�4���z��K�<���.�+|��(�PA�t����	^��a���9���܍�s�����ì$��F&�!:J��&�༥n�������M�n�5i9)|�E�(]��-BG��.�-ԯ�W�+��.��L�������$��;v��14���9,����񠦰v�	�_������wls�	�/ٶ�i��L#If����k�`���
a>�j�TIv�H�]a'��8b7�H�Ə8"�.�0���Cvz������VzϧGOL g�J	q�B�n�k�Ym�Rf���C1lm;�=L�#�LXQ�V�2ΕH"�G���MN�|�c��v�"M`
m��04��7�ى�$ؽH�A�\���sm�*�!'�#-�9N����Ka�j��q�M+ ��iA��,��)fn�_��;��th�+�ۙ���Ѹ��ci�k|���������ߕ�:Q�5A��q<F��-i�o*��GW�`�������e(D�GM@�C��H�p���.���XA�U��ǀ�n��	�O��$V����<uZ�u�S�P=
}BƢO�*��4���;"�����!JS�Fm�"���>��I:���m���z�EZ��A>;�Q�Л�4�"+��hR����͉ܺ\�HP�̬&P�1j��;bԖ�w�Tz���p���m1T����B��]�W��ˬ�a���Dx �JsԵz��d�M�@)ꃗ����:�H���L�\�1�-�L�9�a���nIa��9�X7���i�a(A�J0�F�zX���+L��'�����
�����Y�I�p�����Q�b�����8��l{0��>�'��B�2�8S��0�������	�s�m�>m�2��&f�i���˭�2�P�03C��b���p���k�E�h��)��!�C�����q���e�\~�eH�ՠX��:������yTO�
e�]!e��d,�s�ZxH2c�X�'�5d�!D�3E��T�b�W���F�vG	Th��c��'�]d�5x��eA<+I�9zVG���rz��$��8,8.¨���yHG�-z�4>�L�{�Z��^��U&U6��=������b�	�;fZ�?�_����v���6���h��z��y�P4[�E���������޷�(��QD.����d�c8^a`˼^�~���n#(��$55R��]G�&��3��W��w��B�;u�_p26�'�~dɖђ�� a��&��=�YaZ��
h�Ks���E�4xYM4n�+s{�،��x�� Տ�ƶ�B2�j�h��խ���)�W�����ȱT�f]���ہc��
�l��L)��u����{i݇l�\��:���\q��	����yo�L���y�D2����j�����=�V�k[�{y`|��Sc4�<�)�N9��,֡��	wl:��m�6��.o<Bt�i��<�Bș�K�;��<B�3 @����pdܘ�0�+�Z�WjK��TC��WdĨiG��*���ƦgG�0��G���B0�������3���_DM�dD����
j
�p=��T�0��k:M��iw9�ׯ�>ø�I��/�(���qڭWǺAUIu��Q�RU5��<lXt���5�M�`ֿG�*�BL�	*։�2�5�oא��9��U�utm�z�k�)�.J��l���ޡ����.�g� ���kh(��[k�@�[]�vi"	�pc�4��&ψ��ɤGc��K"����\���:���)�v�;�����7�1�'a�7
Gv��
!*	&�����?Ul��a���_�9�9���<���]�4�Uc���3@���:(��J�{aj������FM���5���uS�-oْ.���o|��$�(]��nCk����Ҏ\���dx������ :��Y�R���B�rU��`�#��@���)C��B�mۀi�����#��}��r������]V����]z����h���G���r3k-���	��G""7v`�P*kEl�f����GE�0C�8@�����}9ާ�G�f���x� ���� ��8h#��m��V�C�V�'�3Y�`&�'��`K;�4u�8�~I?=��}
�����mb'X�+��Ym�T��g���b����r}~��2�ӳ{-��+�0��ħ�~~�m�!�,A��f�yu��8"꟏v��+л�Y�����E��Y���6�e��9?�\����Ե:�P2�OZn��䲠��I.G�C��c��bV�V��u9˨�N [�;v�GLx��c�f�a��K�)���zC����Sr�Q	`�+�"�/��8[�M9~@�,t���6}���k~G*���4����X���g����m�#O���� L�� ��T���l&���褷�8�Uc��'��2;�`������_����3��V�[�^we2e�ը���z�M>L�Z]�����f���Em_
��7���l�P`�t��-���`�܋���h	`���?�ܙ���5ѿ&>����زl�CY�E�T���ʢB\�3ƄX_8�1ac�ő�0}��B?���rޏ�v�mBT��gןmH��;�Ujln�X3�+�.Д�]�(�h����ܮ��B���OC��Y9N6(=��S>/իr���\WL���0.�$��
D���'6�r	T��8��"�:͟� Ԟ�ba�u8]%Uس��y��b�9�ܺ�k[��a4 5��.�������<�ou����|+ h��n���6u
��c3-��t{�K���1�����Y��v��lq�ͅ�-��/	Ry�@����[�1PK�>�7D9]���6bqs�^��Y�[L�k��Կ�~ƏMk�uu�kC[�� :U.r����g��W,����@���t��\�"|�=.�����^(�%{�"R����h��#c��6WV�c�����w�E�*���fsk��/�98�</�R��:~����"Pş��ɛ3v�<���C[�����My����e7&�nˋ�v�*z�nc�s�3��Q��-l��~�; �R�Ư�z����O_��Z�{���f���7�����)kMv�-��T����T�}�+|j˥ =i��Xs��$��z�#�����B�|M�t�N}���n/�LZ�䪏���O������B�}-����r�@'�U<����2�n���h�ϫ,�f�^i�V���,�od���T<})��H-����-5L~��F�)��ZM��}���ʸ"� �[+^o���!Q�j��Ğ�7qF�j]�W��f��J]xJ��'�S#N$j�6�{O"I$�����]�</oy���ޖJ,��щrn�رp��4���W�@*gsq�����u�{�^3�(^6|�.���O�֥"�\��ZtwJ	�����I"�]A�$mʋH���M�SµbZ��/��%���2灧X K��-g��-7(NMuu�vةo1�ɧ�)�/z�'x�G�+�b�(��?A�0�J�4�{�����8������GE��_9�B�ObٺSe��J�~)�u-�Zi���Cc�ĵ!�����;^�AcYHw�wr���4{���]L�&}\
�Q�JG�Z��z���yȯq���\��#������AwÉ/[�o%C��.î��8/<lV:� x|���41Un��3v֓�N��F|ao_0|�j"0{c
W̶�\8>a>�����Pcò�o(�P�$�vqyTPAC�_b8�`���Fe���T��,#+��`��k��u� 4#Lu�'�Ms�q�ݺ�b� �r�s�=���U��d8��q�%�� ͥ 8X�jj��!���I��Nm;
����)$2�R_����/�y�5��:7a;�K_��.ʁ+h3�k�t0�aўed��2���:��`)���2Aɍp�t�6,e��E�[[�׊���+6����!\�uWV7	���J�/��G��f�[�1Ǳ�+z��K���Ө���:5rw;�v��Ud{�ѐ����iZ�^�ɞ�l!�7�s�`�1T����4uK$�C_�H�o0�K��7s��[r��$Z�LA���DN����X��죞G Nõ?��:bR��U����T�i�c�toM��GE&���лH�{�eP�DA�裼���$;h�M?d����n�#��8��89�h�SEb4&'�t7�ŷ4My����c�Ec[�YK�����b~p���yw����3YF���Y�)BY�����K(�Hb���q-z�]=��{�F3J{�)NɋeK��Tw��% �f�|i�ë��s�'��FL��Q���w4Z(�G[�g���V׊��mW��%�2��0� �30f$-`Y{$%���.��VF��.���P�	��9Lfz��~������	eƩA9�%�r�����a�è����0eb"�+H��#Cl�"ـ>��a).�>T��
2�q��蝽�kUg�q_y����x�]v|=O��P\�QEY�#�+U(�..*�% ���]�3�]X)��;� ����M�9�P����zO�n�sH�*1;���D`/�Nfy�X��
(C4Ե����$��6�&^���^#:D����u��Ww(��f��R�(�$�9��|�����~�N�G�dB�0�
N/�r��)�M���^՘M�Ө���3�K������G�lmq��*��ý�b]�e��~��8y8�Z��k4ǐ�b/T���e��.R��k,�L$wZ*��B?����3bb�NZE����ڋ�х���ʙ�#_�T(���u;��
���l�6'�]�d�O�{2N�U�J����O����&�`��U�3�W����i��@��7d�WjFY�1���'���(�5e�;?��w���J����!�*�Kæ�#�OEV$;<�ٗ�9�2=�2t�-���
6����F'U�C�fgj�C	q�ۗX��b���\��Z��t�m���d]
p�i��kjbg������@-T`�]F`�vt���@ss�f�q��7�+��t�T�u����|�Ol�ܑ��j�c�  �xrS�O�b���y M���{�M�GvAR�ս��(R#�-;���t�.��X��@�Әί�Zt)�z<�����E��&?�"M����oY��_8쿺?�:]m���
���{��"	����wbU�z�~��B9��EQ�Kd�VwNӞ���*��Z/��)V.XBpJb�?��֟;;H��A�?��] �gj���Ξ6Taȼ��T��j[��ӝ%lx3<�9��6��f'�[��mJ���PS�c�OKWw��JR�g�>�׆�Q���M�����'��l0g�e �݁N�P}��c�\�WM�ْy��n6Z�G�!=�ў�^�;#\o�\��� �ofv������OA��}����>F�	@Y�9/��`�n�'�m��`�垓��[H��R��7�r�x
|tI�@~0���A��!w�c�hc�*�<�-!�/.SI��±�w3A�g-�[��֔��Hy��L)�ϳc.�i練x�ڼ'��<�Ƴ0�	��j0 `޳`��^�[�$9������K�(�f�&��!�}�/o_����W�3�u?HPs��J���vA�d�����p�ȆS�)�]ӆ�7hIw��O'J�����D ��^n}ա_d���� �T��,]N
S��3��K��5�AK>K�NG���+[��$����zK"��|5BBkd��as��2�q( _�ٻ�N��p!�-7�+�D��{�g���gi*����Λ�"�7l@��+��������Ls�o��vԏ�c�#�%Q:A����m���--Z���W���;)�,��Y�JQ��M��YR���EG�R=��4��������Ro����&��|�Ý��l�y���d����$N�c�x|�#UjrX����:������6���6Wy������lP�>�������%�d�BV
7��7`K��3I(�>�u�[isE��1�k�X@�è��4��v.��Z�y+���]�N ��ާ��R?\z_��@^��E��!>�SR2	�y���r
&ET��L|(�k�����L�;�]�y߻�H{�+�6�j$n�׃����l9'0Yp�m�6��$_�Q�w���;�t�.L���f�S|%%�HE�A�V[��INT�À^�k?@���:�>vxLM	�/�v�l<�1NZ-�f��h�Kp��`4��%�<��F�O��"d��v$:�nN�����گ�Ŝ�]�pO�X�!&٨,Kf�9��.~�2��''��(��z����#ʏ70m�����,'x|H���)S0���tʰ/Ҙ��Vت��&��"M�6H�)V�u�� �
w��PQg���s�il!� �Ǡ�Q,b䦆�HG�O�`�!a�7�& ��F>y]ρ���J.F�9���?����.bw(<����o*Mp|kAhb������9��*Ty?�3�)��ԯ[e�~c�pl�~�^�� �],�� �X�|�2atKG�Z]̟��)�c�lbM���4�zF%x'E��v;SH
�LڏQ%�Q��>m�Y(���B�P�m�8w\����^�ҝt�����E����?%�
U]��eJa?c�{.X�ڒ.�Jt�֮D��P�������aӗ6�E��P���~	9羙n������_~�yaE��l#��Uv�Q<VD��DF>Cn�@�~���^�$�����θ�Q��Ɛ�[��r>���v�H���x�HX�q��������[�"�14uUN���'��:Itǵ�H�g���_�������������R\{�'.]� �Yb��T���Ya)�W)�q����I�M�ͮ��= {���JpHF��KA��巵�Fp�Bi��Z�Z#B�?�����
���-�={�c [���˨w��h:�|
�|�|J�M�p�ؔ���s$@��!8`�˘`�G�Mei��hc�H�e�=I��_�n	��}j�Է7��q�g^h)j�z��e�8BH�c�RLM�`	�z�C}f����(�#�R�3��%ݍ�3�����D�5r���*�����B91��=��ջ�z�b���|�-W�e�}�0BV{~��P��l���W��b���J���)�N���5�L�(�6���P���/z�����r5Wx�Τ�E�.8튢��o��}��[A�[#[�>���I������6���Eu{����4 �s��\2���q�l�r�\�J�6���}sȍ��$a��]���U"���mg��M`�Qs=���.(��~�̌EW�����8�����O�3id,���L��Yq�!�	6$�f����dE�6$��(�`���r'lğz���&��f�]����W�O3��'|ʞ2��m��`l���}�TUx��'�Pz�x�a�@�����]��ޯ��SD�W�8��=�؁V��Y���0|����P��e���L�'4G1�E��k��X�rbaԨ��"�5�˾�Hm��@�����3��tZkf�] X=���M�� �P	���=�zt�X�V&%��Ll��8˭�X�A4ZShV�PW=�-���<��d�3��otT�8���eI!U$�]���Z�ꊔ�}?R�g<��@�����"�n�<W3k�Ϩ5H�N��;�]o����|�,l�� ]s���S�Y��R�K��2x<���x��8�֪޿�Ȕ����Jο��9[0OC��/���_�4SQ�UO�d��D�䤶���:ؿuR�}fE(s�KdJ���C��K��O Q I�Ҵq+����p�e�������y�}_#9�mk����2�$�������[/�`���l'��q�N#A��>��:�u �v�!פ�e��������u� �)��Cy�����.;z��wߠF%�-+�*� ���
��t�~�x@�o���*T3?3��D���\=X01�"�!�eg�b�\>n���dc�0o�B�\�ڟ�����c�н4�~*�Vx�G�H�����X�v`���Z�e>s�P���+g�Enz��Q� ���-K?k G���^t��&&�'N-bM*�_⇜��W�Ak��@��0�=^p��@E�An�����bRjurj�B}��Ҧ��m'�5MzJ�Ӓ�����Tq�K]�[O�2 [���t��_�kDS�M�/v�Vex����gp�-���a����O0���T�$?.X���x�����{��
�Qv�O�׍7;���9Bϗ���u�8B?��2��A���t!����HI���ˌ��Xl�	��;Oy?��.fn0�Z��j���4�1]�^�~�b,L���U��������ٽ�74�\��BB�2��~皝�D���n瀗��H:�/$�N�暴f�n��ҟ;{���.s;���+΂�5M{j|���ً�yS��~M��"�m���1F%��I �W�&�4�]_d���{��]��|U���iNsf�%���O
�_��ޫF5�"Y�D��2�V��u��܋����G9@3�xH� �x�(�������$xC�#�IE���]��j��B��Ӏ�ܗ ��}N���*+{��,� ~l���˽��@���6�_Tm��t�v^�#6=���%�լ�ɚ�Jl�c�0�ܿ��@����k��N�<͡1h-H�ӭ"�g����$1�#�����5XV!TV��V�lc�����'p-k���W�%�j8|�j����l��Bu����w^b�j%���}��r�Q�U�}����U���*����4�b;�+]mG�[K��23��k�T6\˕�GԲ������t��]׎��?ź�q��:�r"D�����Q�OH��-����}��K��E@n�� �"vQ�nV����g?��(C�9�j�D#R��C��Ꮙ�9�e|?3ƽź���(?{�ΞUZ�3m

�>Iw���3
.���e�(C>h��
⭸�C77l\0��)0�c([���/��$���`�ZcpA��BO��Gf[;4��g<Dd��E�6H؆�L!���%���h�B��2���G����)!��}��y�EE��$�C#����3s����=�E��$gѥR0AgF����S�H*�������{Ə�%��Y�8sw۳ q`]�B��U�b���*��z���lP�2�O���!å��P��2���H�����d҄�j�z��G����'A��ʆ=��ꈐ�%�u&���Z(��ߪ|N�L������n��6�J�ɒ�=�7�����Ja@�-\�e��Pv�G��Ŕ6�s&�O�A���[Ӹ)�M"��s
����@8�6�D��v���hǁ����+�$�����:	,��7�����ĕC�C��/��5���ܳh��j ����y׃��3w��I�`�FKۣ�b����h��J�a���R���z�����V� ���������7���q�ĥVD�QL�{{�񵘂dJ�^e�Mä�TY_�G��x�����fq�)���1�
��6I�0ؠn�B
"���*�#������(�4�4��iC�sNt�����h��j\*���
��j-��Uޒ]r�I�y�N-��s������qTJt�@�ƃm�e�� t=n^��DcŇ�`.35��M�C!C�SemW���$����߿/�������:�w�I�5S3Mj�	��{���ɹ��F@߸��SGn�4w U�S	�Y:�āZ��Wļ��1�hW,o�mI�/��|�.����c���}r���P�S����3ߘKrmM9=�44xΔ���;|+���8j\��` U�S,��8ȵ(��)��Aă=�kr)�,��qQK��ٍo}�ׂ���Xݼܠ�����u'����#�=�r��[�s1h�s��,�4
���#��.�v� �[�uS̅��F�6���g���*FfK�ko��dp|���.���Ev�ʹZ��f�hq�>���-�����g�����7�w�	�.'�1h����4X�뜦�u���W��pwg���htи����3��y]hi���2eY_I��s"_�:@��������Nj���X�R����.?�p��|�7EMf�������u���|�Dۻ1�) ؛7��&��Wh9�g�M��^�3���$���DڡL
�<v����,ݛ^6���}r���q�{-ו6*+�{�ؕ
�yv�)�&E�kC`b����;�ao�&z% ��Ṃ���\�|�8,��3��-�\�1D���@�����|�{B4���'���&+�J���Ut"�T���J.<f&&�0M��hp)T�$�y���y���@�/+�X�,-���$�o�j�����{�zy�TyOW/�\a����L����z0��~��P*0��r��,������xXD!���:���V��W�|$HJ��mv`Em�J`��� ���v z�����ަ�����:��вv��Mq`f{��x��M���ԭe����u�o�K$�0����\�R�aj�д�z{�LC�q����$����O�}���4�>�%�蛝+���*ʷ���05�.ި���,C����h.�S�c�2O�k V��c��;6r%���2��R�>�� 4u�VҚE��D���J����͇��^@{�5�o�?�eWb�h'H������%���t��lwH#�P�U����)KsɎO|��p��K��O�zeMM�<}s0r���lds�7 �7��`ݒS�� _	�'��|;NC`E (�՟�HTg��P��d�R�_;L�6�^�D�$��}�^��|\L:Č����a���.u�!s�ص6n��>(i���&cƖWTg2(�Z���}ګ7�<���H*����m�g�^�@��*�7�q@�L�5r��dIw�[���̵=?�<N�Q�`J_��OЁY\���Iv��K�^����~pe��u_�.�!��R����Ld�~��;�^`6��O��i��g4ñȮI�~&ݮ�$��m �M��o��x�Cem���@i��&l{�+�Ƌh����q��ܦܡ��яx`�����	S6���FK4��8�:���c��4��;��Zγ�u��5׃�O�xϓ�c%KKf�2��.�8U�,����P�$��L��fIV���©-�T#�D�i��� P��ĉ�,�F&�M;n�X����P��^K�h���R��ѐ�����19t�Ď����L~S!��"1x疍K�
�Gu����7�>�Ƽ������.��:�����z�c��K��%�괮���-���>�ד3m;a@�O�!��*w���	���a`N9��f�y�-r��~Qh�&9bz+�o':lyD8�~ߤC⍬�)(��"]O���T������Ϝ.�Rt��@k�[��7�"la�]��I|'����Po[/��qiӸ�3����3�Rs���WN��-�H��n|mo�#���S���-9��z��wz� ޱF��Zdoϧ�Y\ݞ.D�R����K����W�?��f��&��t�Ͱc�S3
-t��%ǖv��jd^M�E��us�~� �mR���|-�~ĥPi�8�s���4�B����-0A5!���5i2���W-����Xd۪�O5��,��)! �a��ʦ�AcTXZb�P��n@��)����SY��{�H)H,���@���Af_=����m�{�S�S�)��'O�[uΦ�	�0� W�-i���ћ�ѷ��KqZ��mM55���ZB�2C��{L�&/Ftt��s�-����.�v��n�	Z�s�Cr�\v�KhS�ev��F��S"!�婄Xڠ�v���Z	'�{�7ן6.��>�I$.$����]��_�)���4(��#m0lS�$�q.��wڢWV�|�t0��\iE!.���Z���-�G�rE�{��y!QC�;5JO�hI�]j�%?囡#V`)ޛ��ǡqC��3U&��5/P���*��$��ҳ�U�>{s�n0�����Hk��P~_����-� ��=�X�W�Ϭ�t�ENxL���oA�'�Lsh8���r�����������k�n�l/�_��*��j"D}^��_t��^����y�R�x��������6.s k���d�o�����d*-X�o gs�^{rC$?壄������9$�[��~6,2��C���/�`��e���\Y9E��L��_^(<C��B�����b�p����Dl8��F��ƚ���X]$+c�v���@r�K�3+���jC�:��q��<Y�F�u�V���p��=-X9ZS^v�"<	�fy�GEκFH�+�Bee�1�Z�JA��~�G�%=_s�>x��BeCI*���	Y9���=`����q[ ��������.����~�|���������ℨ3jRD�i����+S�o�c����N�!O�!!_�����z�Rf	�ՙ���E�X;�����/DI�Yj�Ѐ����g��\�H����
R�Y���כaRa�*�զ���ʋ���W� ����Ǽ��D��ù�vɩ*������n��w̳���ǌ�U����ɨ�F3'+\ZՐD��@���m���y��,�`��ѣ�E�iYݿ@?s9��0-�Q�x�FV`���<�iJ����`��h�1Ed!y�W�b����� �T.q7}ơ	���_/ %7v�Q_��ryp�YT�t\$����?l�5�/��x���ԅ�{u�؈x����X�C�	7��mw�<��U�B[Yn\���6��Q�tA�i�{���In��q�u�g��ƉS���.I��@#ͫ���4Z`-���He<����t�*��Kì[,�JI6WI��ۤ�rqw?w��5\�T5����$�|� ��u}�zm�����=�v2�:Q�I�U*a�m
U��@��̎��Ԗ�f��hfBC��] V�(1ǟ��E��3O�2,�~���瞝�ZLK֓ ����f����IT�-2���<A5��(�K	��\��}L��6�_�TX�-�����rbE/�������!���F?�����ȢV{�H���8�4NU�Sڳ���M/��@��S�e�/3��|2v�@���%�Q�Ɨr�%��u[��H���i)��0���2=�6J���,i�6�g�nd�8XY~���\:�p�>�u�{\8��}ڨ����D[���r��b��w��k���j^cg�t{T�*]^��?y�N��oFܩ-�H�JQ�3�
2`�!m:9l��k2�߫=ܬ�=Ap�� ��a�n92;��&\t�k1��lg4�j���zP(~�0�)�ɑ�B�ťT�-&���K7Q0;�3!����w�`��L�������ı$�+"���z���O\�s��Ͱ�j��4��)���H�A���4u�^鯓mp�q%�H�T�~h)=��Y|��5�t�_�����")wP�]1��u���1ϲ��p<*����G�,���R����J�����R��S�dʮEʌ�"]�'j7[e0\r�QD��ⲁ���\S�����+�ВcR�~�bˤ)DFБ)y����&�,�T0w+�ĿU�t�S�IA����)BGirmg���x�}~-��]B�A��g�+�${�}�S�Ad�؎q�q�����QB��qQ�V��8~@+W������^}�o�Y)[���]�0n>O�c.Tf�h�z�s�a\������M����~�����DV5�F�_��S����(>��[^��L
�5�ͺ�k���'73�0j���O��ӿ��":�R
f��$���<�(�Z��][�+���������c�D���$K���M��жR������ۉq{�g/��)�$��͸m�����J/;���ϴ�v�O+>p�&l�0z���3���q�"�^�JD��E:�$��
v=��6�{Ю+H��j�=�.���<�C�O�q)�ҎX3W���/�����_�Q�	�S�|��9��R�IZ���P)���?#IV"a�?RP�Ɂ�1�T���1���dC��)Y���d��3��s�bɴ�5ٜc�=� �/Ud�S\/�Q�2|���Ҕ��)���X
��R���K
��f�&�������.�����t��M�cݙ0�)
L�e�?-�M��k��W�-"�<$[���z��!M�`�ٺ���Ŏ�Up9�c0-��!�c��̱��J��+7?e�t���Cs�s��q��(?����hz��A��!Z|f��U�DCXf��6��8�p���^�U��~��b�˚�f�Ǯ+_d����>��f) ]5Ϟy��_����38G���xA�&�A�5	���=���"����5�LF��1����!�\)�&����˪a)4QFJN-殪2	J�bz�Rr���� D[�t�ǿ	��Ǡ��ɐ3R�Z;Z���*q-���.[��Vb�+F����\l��W��F�>�L�J�֟�Z�-��7v"�Q?��Y1�C�12��ԯ��b�{��j�䥎�֞���5��\�%?�!��m(b<�x]z��^LR_���꧰Pq�-��X쓙�O�N��KA�
��7R���령{�h朁c�,�C�E΃��)�m�;�r��(1B�b�,@��dpnA��([2��ǡ^]9������5k��|L5T鋡�jcz
�^"1�/�����	��|�4��C�aUd!2�A�g�kdEG���Kq$p����P�X���KĤ�E��'�d�\�������tϟxo��&��_����aQv�֜�Ndw�	!i��ä~�Z�F �����3]x�,�fze�������	j,Ŗ�r���� F���YS��"��.9���j�a�|9�׹)�4Ԡ����ϳ�����'�,^M�f��-��>�������BLJ�� �*p(�֕U��
�`��R��ys[�IG�V�fkP�Ɩ/���v�-�ir?KEKoKP�o<˙�֣�~���긑�%���4�H�6<�R��z�9�ʩ#�Ӡ�| �FB3DO�&���4�����ǭ0�.�gi?f�qA׳��xMʅq��TE!�c�O0��c$�kcNڇ��#�e���O(�`�Ó)m�BG���4}bS܍�b�"Z���5�0��0�k����0���P���n��ݎg��:TT[�����A ����d�>alU2%��r)��A	�Ł�1����fV&Q���n�N(s�893���a���-k[o{���0�JS0+�~�wnf�f��h��M�'����D�;�RߘWq�ZV�A�p�����u��Q���j��u�@�����[��V�=j"�+�vK�J����\�o�8�5: �|ԕc�C.�-"�5I$+����T29�u��|���R�<��L^b���8�b��5ys�ddyL2x},ׄ�s��/ހQ�0ѕ?��	g/����yߺ��\8���d���-Ꜹ4�/��s}���W3�Bn���g#�#Ix����)�[�s�qB���~Do'u3ޕ�1C�O�d��!K����?+ �|�V�O��o�f��#iI�pk(�DM�v�-5$�V����OqPn�u�?T�W�$�����G��HC�q���A**$d3Ļ�h��!�U�ޕ���x����� 8�� ��K���߷xi{R�,Ds�O�Kj��W�������0�
��Ѕ���yRs�cZ{D��"�^Xt���ɱH!
�
E�E�׿	t;���q�Z��m�}��.*,�z34��)|h��h"����E��4i3Vm�z&!i���J/ ��,)����Ҧ��Yls�-;J�ؾБB�9Rz�I2��T�if�n�h��F$-|��z'(~���=h��/"�!�NC`i�Q�8���aDE^�K�������bj���v�uW�Ὃ�,��+G���^�u�&�D�Ԅ�T��£LB�ŋPe�W�*\2E4��bYL�G��������d KQ�'�6|�t���p�M��~�!��HJ��>��C�٣�5 t�Cu,։^˼6���P��G�s�*�!��,��D�}��G�5S��}>�O1`TBږ���m�琣�`9ٶlo�M����x�b5x݃7Gv)�d,����kІ��wQb�]��(2$\��׈wV��f�U~�#��݉�-=r`-��A�.P�?�|�LW{L�\\�;I�����b>�ҭ#�Z|wNR0il�� ��\r��q'օ`q}�bo��]�X��U�([�cǃ�N�Ҏl!F����Kp$�Q�_@R�(���%Ƚ��@$����z�%���e�.�(/?
c��Mt���G*8
m�d>��������CU#��ܲ
)���?�;)Á����Hg��!�	%!e��d�h����#��*��f�C�X��.�9�߹�e�w�n��ɡ��C"�����{U��6�������&��t<�����W�U��%�O6��0��%"_[1J��l6�fφ���Q�|�m� �<[d{�=1�Fչ���d��Ǡ�EɗA���)�F��ι >�,��_�?l�/�Z���u�.�JT*Zv���lt\g��d(47�(Բ���扑�P��Ԅ���㉓l1��-{�lkp�ă�l�����%�DQR�A�j<���x:Sm�J�֬����,���n�~���(�}�3�S�wq"����m����yR��,�_Q+���ǫ�UE���*|J���A�׀+k�{VF|}�4���Y�t�e���D�ucK�ө:-��,~������pH*��T������, ����Y�t"!L���G|[���R�d��Po]46Hc��������������&]tK��R�L�Z3���x�si�~R��G�����e�@/�Z�J���ɞ��;�"�`���0��h>�|6�]%�ܴ��ɜ�]����>��{� ����,�8ZU�}eCw2����t�8�9��.��A����k3VS&���ƥ�����ـ\�z� ����!T��N!���C.`�y��({�E�R{���<��2\iH겖�|��ߕ��Ţ�C�m&�x��qkF��Ԗ�6�"o��d���AS=��uva�W���X�@�Ny�3C��"�	҇ڼT�1#:>�k��-��;(-�a
wK4�[�����m��;�nw�ٲc�iq�P����U&�㠳3��J�{����V���05
M��m���kn+r�d��.5k1�//,:�c(�\�cػ)>i����e�R�'JH� �G6J
z-���&�86b6(���!E���qb)8C�;��`�*��X*�j:��k �����`�0K��*	K; ח�K�ضԝ!�++��Q�$o63�>ș����,4�Y��{Qy���!͞E��d��-��%�_q�S��u�㟠��,G*�u���`�b7������S{k�`�Ig�/��`�rӐ^�����Op?���F��t�3xy�Q�y�g�k�[��>�����,�MFuʻ!'���L5��?Uc���L�-��Њ��@�En��tt�h�>���6T��d�~ �˖.�#B��B4}�*Ԙ�tx� �qh*�V2Nb1��&$��,�T��1��O���;3VxY�({��/9�G��>�@N9�L�׶�/R'�T��͝�Q�Ug�t-�.aR�\�L�K�z�@^i�o�&�����#E�B�Q������-�禥{7zshQuB�:�;�
Qɽΰ�G9���"̯I�4Q��G\?��u+,���<˵������ir�����KS��'u�5s�Pw��^m3��nXf@������G���v��<D0֔)��];�}�|�D�������_sqN�q���{�&Q]����I��sG7��4��8�T�3#�8SguzRrv;���*ǳ��B�����Ëϰ*|����t���s)��.p��*=�#��Vz���3��Jvj���V����d�34�!�|N��L
�������bν�cu��/�/SPt���SA:��`�,b"�n�����q�@������@�����d��*�%<�)��u�Ag�\��cBK�$:~ǯ����Sp�B�mP��w�贊d/p��4ĩ
Z#��U���2�5%�#�Ɩ�0���R���]����Nʌ۷8,��D�;p��4sx$�_��+B E|���M��I�S w�s>O1���e���C��i����d�s�MPT<���t"g�� ���zl�;�2��Nޖ��WC+��e!����i���U�	ȕa��@ղǠz��w]=���m7���v�vE�S]w�H�= Z�Ml�,NS���>mG�*L�-\(]�d�%m�ϥl*H�H��~�4y���2R�{y�$�J �jΫoMk�^	��]�^�r�9��=�J���S4�s��B�	5V��d���[JD:��  ���bG��^��B}��\PR�Z���	�ٕjf�&a���o]�k���w�zx@@a�vqzK�2�l�_����x$݆�uF�&!0�7��p�E6����2����I]���ULWiZ�{>r��;14�n«�^xl.~C�3c�HNJ>������z��GX��.�1������S��h��))�r���;.�-=��5n�	���Ӵ��g�$��Ď���ӷ�w�w�K�cfd���e��?��1���xH.yw��
Q�� �}0�Θ?���,��z~��QJ$�������l��8��!*~|��g~�'H�s���#P�ms�t G/D���&��p�s�7�=�Ǉf�<�M��w�!Y���ā���r|]3�����(�x�AƸ����ů|�M@�����L��s.H%�!�f�(Y� ૡ-����`�o_ν��,
L�^�B3�2�@�ͱE @��z0F�,�\�����uj���E{.6X��!$�:��9
g\��{LI*�T��-�#���2����f<锍i{�FH���j�DX��A5����P�BR�.����4���l�^�6�^h@���/n� t�Ɠz���l����؉d=A�|\�Ag[�<��$�1�P����W�.�j���T�(r��q��7�	��*��h����֙�~���)��:�vi�]k�>��[
�k������fʧ�����U$�r�_�Q9���%n���_���?�{�T��K���o�CiC���b�
��b*�j�,�!L+q����c�~�ؘ]�.I�����F-Y�{:	!���c�'�=���-,l��`hf@/�d!�P���|����f��B_���7u�Mz���M�VV]��.�9ttA�6=������]_�\v�㎉a ���n�9��O�a��d�[�e[� Us�) 5��z����P��E�T.�L��<7��Ǥ����h�J�R�=��oF��7�h��F�8�7J[�ɵ�U�F�Ҭ����.��Lt�p#��Y��?�!�8�vof~y�T1]^I�Ra��v[�]J��ڼ*ugS8��U'�F}�]���G5�}Aj�\�E����L�O�u�h|K��}�S䏜���GHhN9�oA���1�y��6�(v-÷H�@���A�cx�'K
���d� oý��)5�N�x�|�������u���G���K�d�b�~�"���Pu]`�
z�SV��T�k��shm]���|�&�|�ʰN�M�.��БWjF�0骙�-8�a��X�s�I���N%�?��������8̕y�U�m�W����*����]P7.�9�4�MQ�o��m�с���^r�bn�?��H�d��B������/��0܏C*�bӛ)� >������FAom;�'�~�aěY@O u���M}�dw����A��ʁ��P��5�], ����`q��Q���������x�G����Z�e�̄ă��A=��&�u[4�I��NL����fxb���e�;cΕ��.k�3u��їR�;�ŕ4ѽ�v�7��خ��e`O�+4���S��V}7q��z~���T��
�	�� 0���Ty��m� �UHy�p�� =���|�����K��٠/�WS�BL�T���g������kB07����W�d�~;��D�XXd9Ex�V��Q���k:d"�.�~Y�ֹ"	ȷ7�ӄ���?�f�̪��<�����2Q_��¦ᡦ6}h���" �wo���~��w�6���<b$��B)�������!ϡ:J|
���(���������I�?�o�X���w^�m���K��)n�,�E�2o�&%qB��(��ϗ�?8YY���hR�w�+E�j���X�V�|'���J˶r{M���Et�n�����`�,�#�H�2����']&i�@�wTd�"S	f�XO�ܹ�+�"aC	���sP�����Ù?!��h�@%���ߝ3�
���q�C2*a8*}�Mz �eJă��4U�̉DZe���>W���ոQ���HwmK�4T7B�@��`\��Ҵ6�rk@�`>����<�$�r`=<ͿVR�W5���sϐ����YB񾉀��5
(���������W��n�%�%)΋^L�r]F��?69��$C�����.J�����u�3�-�/Z�~���0�,U�XL!��FdgV ��?�C��������7`��h���:�Vq�?�ʍ4�r��a@�ݟW�Z�KE������k�R���%&K'b��nvG���#�3;�zGr�n�]���~�%��.I/�M`pX��LܲJ�2S�ނ[�#\�,���%",f�xҀFЦS�?�$Ɣ�!nm��^e�/������=�j�xF�YԾ.�A[�Zaf���Ut��S��ƀ��x�T��mI��o�<nR����Ĺ��N���ht(��x����p
��us���?O�͸ǀ�)��	iQC#3��-kw1�އR��_<ί�0�h/h,l�Ku$�M�]��6���##S1pZ�{�M	�^X�R�����qFZ��D�`��8v��������$`�'���)ާ&/����c�[���阹N*�	��Յ�!�o֬�		��Mˇ���r�e~��a�Qd��7����Ю��,]�%�e����7�8&wO��G=":H�[�Z�s}o(-I��X����"�m����t�w�X��,�;�-����P;��:�T������Pՠ������_�=Ib�W�+*Ί�X������{f��O����	�؀r8��z;{��$D��&Cg[�Eqd
�e��NŢ��\#i,Y�X]��#y�=��8��K��ŕ������{�X+�
Y����{i}�K8�V8j2��ƹH����x˰�6�UC���J�\�EM�O���_���0�۰d�f�fh�$�0��BF��Nr��WG�ru�I�#�{�v��<r1'�^�bQ�����<Ո�9=��)�Z,��{]ډ�.����8������qi6n�F'��CNd���"��GV��c���:�R��pgq�UjR�;O�B';]��Q���\"��������|�o�A�=�}��vf4�GstM�Zkk=�l�i�?��� ���U�FH�	��>ݑ^~�n���:�ɲ�f�%hh�N�F6X��*5��%2Y4].�^���p%��z�eyĕ����}	�Z�L�	��e}������@��u�4����?b*���
�0��%7���/x;��7���1���u��05����--���Q&MZ~ ��.��*�t3��z%l�}Ԋ�u�8�U��������u?�>呭���=8�P?᷃ɯ����u�fM�p�D཯�:�V�hP���`@�
 �+����B�֮���1A]7�7�(Љnd9�A&�'�����%�@&_���UidC�o��$����������{S��RO�Ll�lm�H���s�6K�j�[�����qᖹzm�S��6�a��jJ����<耂UhVm�B�Z�/����_57�l_qB��#�DЈ�rqQ��(��O���Yb=p3���b�t����|#�2����Ea�F�M���@�9���/������Q�~�����\��UyZ�-pA0�)X�N@����tHR���yuv�GDE�t3�ÞI%8�*[HݾᇓB]�x�Ѿ`v�ǉ��Q�K����ȿ%Ă�� �J�$Ư�.=�������4�����]K��W�Fxx�����X�^j�{8+�r��N��8��4o�W����5�9u� T�]���6M���/=���Q$�e�����vp&�/�U�RŰ��t�h�ۂ+C3 ���X�2�tA�'�����l��88������T_�d�,H {�Kh$�z7 *������l:���^�I
��Ȓ��5 ��B�Xs$P%[D�3�@����1uR���e�Yь{�1�ox=}zB$�����B{R��ݳ�荽��ې� �0G�V����O�/��}��R��V�i~n��?ث�R�6��,:41D��Wm_��
@���樣fHhz9��+q��Pt1LD+ѹt����HHo?�@�[YYV��E�����V#z�(4��`G�D�d�+�h��,�N����=%��.��n��L�PA�f����]H�R�P5/d��2z	a�N�A�}�j�A�^�lX�C�}>�a�֯�r}=��҅q�3���7-ܲJ�UX�hh��>�'��P<�<������;5>��(b�gK����(_��tX��m��8w� �����'������lM��Vf�)�E}y�J�q�%��Op�K�=��0@��;͂l��,�"�H�������)���g��'� �<Q��dߌ��!a��#�l¾Pu�0I"�7] 74�������dⰟV��~�\Ti�����`a8�*�t��`��*����|�b�����7[��!�|�/���(�o�1�1E� ;0p���/$�T�m&���6f�X�N+(�iR����$n������V��*��^>;��{j��'��r��ѷݶv�wv:�l!���t�5Pv�� L~ތ�s���q^�MZ`�����ݟ2�'��Z���x(}��LyţG�W�O�2_d|9�����N����nQ��_ˆ�r�d?�+pG�[`��#��w���;�I$/�����z�7�"|��<�/U@�d��w5R��a�c�t߃gӮp�5z@�&��%�^��)\�Q�cf����&䣁�MP��{���	Ƨ���a��=��N��ܖu�y}s?��W[K��B{g ��B��Pν c\����y`>3�iSM,WS}��%L�`Y�O)����Od�dɯ7��%��iGc��>�ۥ`��&���<B�ͲqxH��U~�Ku���5҃@s>�|��3��/?�6oh�����i��l5�F���:���y���3pi˗��z���|JO��x<;�-� Ԝ�]�H�7���iڍn`V[�����H�Y�ĩ��_�8�N���`	z�(Z?��HPj|���x���A%�o�U��ײ�k�)�XgD����]u�$�W����TO�Zk�^b�k��7����/�Æ�ᛰ��@Yב�x�Zw1���$���hlM�Z~�����ż�NO$�T<�*��p�*w��Y �Z�����Ӵ�8��,���4�꯾�q=Zypt�T���j�Jf�}�[��.�uYYb\	h\�
|��G��t&^�ӽ� G}\�pQ��P��������Ez���	-�ꨇ��8�up�V���H�Μ&abx�a�O�{�[�'��<s@�ʯ���wsD_�zY�B+;Q`�UX�ԑ��-���"�<0S�Z_N^V<Mۦ�9���]�<��Z�.���E���NWV�dB�T=��у�rϱ�$�6���#Jq���v�Q��zs�Y�Z�G�Ь�D� �냗��A�XLk+��'}��-�3��4B[R�[��2Nנ��`v��E�'����Vy�d_0�A�a*���1|����J�fZ�1�Y-^�1[��aݍ�){27�t�h�Kc`���U~����K�ӨYI����ڋM�v�ߔ� ���ԃ��W�. :���8��j	��H4%7�3���H)����x�;��h�����\�؅�U��Nh�)�V�	�lY����k\�lc�9��#��Y�WT�&���O/��_�^B!��E`����c����46<Jy��� �p,�����Oө�T��x${i) 
ο�lZ�bU��&���<oƸi�x)��Z_�B�ɽ��^D�SGF�2���)���x��҅�90h��LS%�\�EH��:#��562OTI���@������ۮ��b� �On��}��_�8��X�s�6��^��E��y�+�}��
�g��y4Ŵ[0x��R�(��T��n�dx@��A�-_�������ǯ�z��u���D��.OHN��苽��v~���#D�`_�.F���	8�T����>S�6LJt��<���a[9��t�(��X�a�%	�������hc�����1#��]��z����)/n�,8�?�ZvH�/f��q�m���u�f�|�ے��;aޢ�E5���]�3��$�([�E?��T�N����l���$kc}�r E��?q+i��x���Ϸ�}C\.n�LZ�q�9�"V���l�#��C �jxÿ2�I]��A	���Q}�C��л{Ɯ�vB l��M���I�$Op�;�)��u�YL�D�s*\:����^�k�N����ș��M��U�.�7.�#��@v��=��z�'5�V|K��t��>$���F��I�����,n��d�ﶡe�8�����O�L�ц��4a����w)9K�@��"��F�G�s��$+�s��<�x��=}��~�й�V3�Q����o{.�U�$��F��;܊uiIj�f?�9���V�E�hh��L�N~R*�~�߶fG�=�͘@'꘡�ݯV��?X��X7}�VN��i4��6���j���D�R=�����R�u|�E!�'����d��bT�Ǻ|bN��T�nY���ï�����+әG���m�_W�Vh��[m����_��m��`����Oi�s���;�����yl�e\�9����AӄK]�5Pp �폘O�F5�n*"��I�-�H$'����M7����3�Jw�Z���B�Y�K���|���~��~��r�臝�	�d��M��$����c���O�R���
8/*.uF[��Wә��� ]�:
�̊R��sP��������'�7Q+۶�t�n��t{�:��ɫ�7Kg���4m�2o��\b����	 B'���%Y%�C�9�з�㉨p�v����"u+i��~����̢�va^���Х�'��O�wJ]\v�i#�󕎨:	:�7Cz��I�AlD$t��{��ye��Ϭ��:B�ΝKS�?��+��r�⤳��۲�_����Z����y6I&�hb~P���<!(Me|��²8�d�2^��D&��	+�m�����lԙ��\�$ ^<��<st����&�o�����ګ�{ x�����)1I�Ǘ��|�� f��Vp&>V�����g�ܻҊz\�=El��81�Z`u���7��/�L��+�)�=[[Z�k�Jg���?t�Ɔ�+0p$�jq`��B���Yʱsɣ����Zb���} �#��6�l��	����VÊ�wGj7a`z�����}�+�FR6[>���:p��=/N���T�CD����{8�
�
i
W�Q"�.����r�A��gtP��`��6q��I�CE�cЇ����
=s;�|�Q������	@�e;c���1ɓ�tq��D��E�E`D��#���5�^K]�
�'�5�WV�*��N��-���mq����-�kHI�����u����H���.�B&I��	t��D�уJ�}���[�^�����j�Շ�}�I
ϧㆴY��L���F�IV>>��{�<=�̻A]�84`�����J�~8��/��Q�҉��a�2�|�,���%�|��I;��8����F���h�h�ɬ�b���Z�*��Ec�<M�#�Pv�d�ؼ>m�6�V�l`D�� 90P�Ğ�<���;tWV����w�;���7Ug8�R���!�1'���qN@���X��Α�@�µ\ظ��!D�1\�_hq~�7���1ӏ��ɣ��Y��p.���H�<.�	�Q�5��`?�e/x���_����p	� ��Iy{����
I�+n�/r�}���=���(��:=��Qlq��K��ΦC�����#�٪D��,��?����m����YE������[��	��KN��<g����J&c��O# Rk�p��/��]��Ǚ�Q��0��k:��M{5Tԟ"��T��������i���I(�~�Ɣ0������89�gL-m%�
H��D0�:��9�ܯ�.���'<µ�R`����@��l8�He����'��g�ϲ��&*���i��)�/�"�y�C������C*2E]�}�Ww����	��߬?e�g+C��\-����S�H��䰐^`��Dp�Z
�/~)z����>�5�>,���a�.&������0J�W�ïӌ����*��kh�(W(�fG��][�z�;7|o��6:�������Q�Z�Hx���P��8�+J����$yr�ܮ�ok��+)�PI�v�W���z�0̘��6���:b�����{H^��mm+r�;w����d���YK�w�@���.-9FB*�̻&�ѭi�H%9��<��zP4��S�۞B�~��řܸ�i��~�Kt3�y�'�ͽ{�fȏVͯ\w�.I�E����*d�I�6W8@�.�Wˬ�̫%�ɍ"�������͑�n҈1�i���W�R |��[������-��@����G���.	"�/>��� &UՋ�j��r�� Xa�yqlFL�˧�����٥���Ǵs�7��'���y!���.S�ɂ־c�8��1��mF���ӕiE���I��e}o�~��$Q&{9U�,�����/G�}�7C��=1�:�� F���ԯ/�d�q�8�{�����=�5֔p�N� �y=Y��x�(LF�f츢�=��>9ąQ��{7]?��A&Yڴ��)��Uڿ@/P[�q�����}�c���������� ���ߺ��zк��k�p���8�C�����R��YB`7�%H,&��/��`�����4b:�q�i�<E^F�� ��*qOv>aӐwpE��Ti���F�k1��O^�6�M�O��_>3��L�ȐS��B�jQB�4��Z�sU��3��f/����	����b4����-≮�c�<ZQ�f�/���u�j�tp����Z����mh��8��N�#����G�zcC���E��<^�)�ߠ��`�G�9E4��������)�Q�'��ԜBI���O������ǚ��\�Ύ�J�l�q����PE��e�:��<c��r(�h*�j̡���%[��;��N��l!N_�`3D�.�:�/}�Q�4�z�9T_�󱎘�qs7j�&K9�`tz�}�M�Y�x�<4COX_�ϋ��!	%/f36|�-`6��K�YVbVB�3@�Ce��O!:�ٛqQ��j��7�o��z�F�ng�3��r�L�7�] ��}B&��.$���Z�)`��R��N.Ǹ��zQc��XiL3(v�mc"�1�n)1[);P�0 
�3X _d��J2�� Z�����ʥ`��Ӹs�JA�-����)}Fz���'���?�M�[��d����`�|�7����=%W��*�GELupI�\<M��PM|A������a�i3��$���e �b�������р���go�p�AFtz.�7X�zۓ���,d���L'�u/WA�ry=+���$������8��A�(ؚn/�E����4BI���p��QYS�=����m�_�$�~@k�Eװ�����4:'i��QB�*�8���jh���	W?�|��F�Ro�JV������d+�!.a)V�P��k�ی�/�M������N��ȯS��J{,{�7oх�	^RE�ٗ?��+lE�L�&5&J�ѯ޹�Lk&^[L��=��_"������ ��G�4�Ai�a�7�y�+�;����F0�+�LO��57Kn�U�ڣ�Kd|�3Jg���
����l��ۭ�A�������$�>I� ��OC�اk���DӲa�6�8 !�{�'�r"��B`G".����9\���u���BI�pBPR�|M>-A��4Ѳ\g���U1��})��������A�UL�'�ld��㜐��p�=�S�J��5b�8\�e2�܇�-j���0aZ&�����1��ni��/��3�+_�්��*��@ �mU,y���򺼢����d*tHCYi}k{��$�h��S\)y!�s��g�m̏��9�DC/=8�u'��jt����(G�K-�!qM��_��X;7�p�f��\xI1����� ���}*"O)�X�2�)��`���%���Cp��`i��zj>�zp���sy�V���&K��9�h�[V�p$�G%����X"N"��Щ]bb%���d׍�����!�͵����0��E���pe�$7� �6=��]%
wL��d�t0�C���%����$��K'�f�]�$aٺ��MҤ�X+��ː7L9�S���2�Z)�X����lE���{�����̶V�n�_'v�U=품����mI=RK�"��w+PnX>tQ��T1GOl��g9VŞ�fI�R���|Cj��,������9[��^���+�mx�Z�LMs��'-4�9�?�rڂ�(KOa_��ƦLN�iW�ұ�孰�d7��f�����8��M��O/�L�Y/%�]=㣳ց<a�R	�T�lXTv����{�>[�(:�o,�����l�Һ�kh)؝ Q0e�x�� h@\. HH���,���
���_����z�᥾>7�q/��ǌ~�\�YW�����QV�Ȑ��Pv�����bI�d9N���n�
Ej�C��?�r���ݨg�/�	���W%07mU��	l�����SӫΜLz\m�L��dw0�`�N��6��0o�O�Q���D�wC��y�~�/T;��]��20���l�D��oɲ9Υ��O{����V���W����a��ڛ��Ρ"҇I����I�u�곤"T�����~�Ьv.G����f`�p}��Y���)�p�Xrz�Wb@�?���R�,�ԙ���p�'P"W������+�%bU�0P�K��9{(��!� �b�8j���|��(u`��,��3C��~�Y"���R�+�5������O��V-��U���y
�N%�t�-�;����̒.ި, �������W�q	nQ���@C�D��5�C=�Yd	��n�/���^!��n/�$�v������d2���?Ƀ�g�H�97�@�X��`{/@�W}O�E�;�"U�%pOWب1�����#mS�0���P!��p|o2R3�)n��?�q��,R�'�b�~MK�c��Z�~'XNǕq����H�
��5ݤ�VzUME�m�v���9S1B�6�9�G�a@��h�E�r,�x�2�+<���zCT��VE�j�8JqY7�v��5��9����׹k^r`2����8P�e�bh�~\��e�*Qc�9�w���OL����1k���a������ϔ��>B�7��� 5ez���B�\�'~E|*�X�v��>� g�Q��W�����[�%Y �"s��9�6h1£��Fsx��l_���^;����J���klp�.���+P��s=6��6�h��&�n$J��LH�eLZ7�X�r��kb����<�!�@����:k�z����CB(K��+;R��Z�ׁ!͐l8;Y'�gO�5���s�-�O�u��!��ݒ2������]8t�`�����a�]�������'�=�S�|V�C���/2~�#输�@r��N"�E�r����(I������_�d#dC �@�*f�'���P�[��+'���2��*�|��'�d�m����-m1l��%�g49�X�Q�Rd�K�pM]�D�t������u���:ث�>��'4�����Ɯ�v�Za��]�:+�y��Gn�l�7���S��~�����v7�`�槸"	��Cp�R/�A���&��qF��cf]U ���]��FHCL������{~�R��# �;�C�zmN�>���7�B�2���j��"<�˰���3���o�A��/��?�d��8cz���b�K3D�k-�}S���(9���`ZY���>�R�&r=)��� Y�+"�tc���bZ}.4���"g{bȊ�?�3ӭ�u-��N!��/o>�߭^�0fJŃp:z�'@Jx��"���9.6��-��#�(*6�c����v��CY�jk)�!���o��0z��Sa��� Z����J�qA!B�6&q䂕�%�ڗ�*�G,��w�e�P�Ӥ��.˙��8wO³R��p���h�O���m�
5L���kO��:�i�	6��C4���w:^
��x��ڝw\N�˯&[����!�������!E�`��x��6�M!�F^�+JiWyR��i0�e\{�\l�̢1w!u)e8��0���:��ͮ��uywf��KX���5ڪ���l7���c`d;����F\�VB����cv�V��*ۓϕ	�'��ĥ��3�3�j`v|�o�虮�$�s �����k��\ ��C�dB�9`]5�\~y�/��`> )��v����mrH�^�M��Z�3�1r��d�ŧ7a#��;�����q'�-�P�s�����+�y�߲�������}���̀i�Q��/�[�% V;�[���uXD�4`ͮ�/�v��IT�+�����%�9�3��sd~y�U-��r���VZ�"�Ai9����&�=N��鳣�Q��志Հ3�V'���������:s�f2"��4�ұZ��@���~g��ϟLSY��:�a9�������w�N*354�uW&hۗ{[0�.�6I5|�#[!��2L,����9�8�W�w��w�ZN�b���}���r�A���X��գ��/�$_���t:m��!�������9xj�l\<bE���.����eV��n�kg@�XJ�E�N��q��X�.d��6L^�T�Q��T[>�#��x�`,y��?�(ͺ\��{��s���l[4�6�ʨ����'*SA֩���G��,=�ħ`J#n���u}��f�nFA�ne���)�L�Bs�����j\|���kr����.�+rH���О�̚����_rC�.��Qθ�o��b���nd�����4.���ֳ��/z� Y�yCG�%=<1r���V�G5[�E�%�?IXJ�d����ƅ���7�+�P�C�r��+o���	��V_*�SU��%1"6�}�ӏ��ݼ�ƌ�������"��)rA�v�[w���H0��?5�VAX����tE��`+|���_]4��V۪�/H�����<�������_�4g���O�&�E�E�wR<��5��jz�v��	��%Ξ�����i���B�1D���n�B��ļ���K��v����ҿ_HX��ʭ_X5,�����lMX����X,+�ؿ<	S�D������|o %R/��tS.M�.zY��������3��=?�G���~9����a�X�#�̜�5�Q��M!k4͇*˵�$��1��:%] N� +�C6Ib��Ƚ�H��eA((S F��c��;���k���R���y�p��)���|����������C���f���6�9���j˶y�O:�gX���K;�Z��I��B:��8܄��i�­����iG~��p�&�;��.�5��9X����ۉ�AP����g�ʾ�I4�a����p$�D���W��y�у���C\�eW��rp��1�D���R�LE���wI��P�'�7k,`�|pW���CZ����JT�W8�Wi���6l��vf�`-�Þ��������+���ć.(��f�K�s<ᣀ�4-WB��\�~�A�W�4I�h#NSY��J�\��3������hb\L2�����ڄ1�$69��O�AwlZ�3��v��a�Z�QNyL�U���4��!+�å'��G��g�dݾ��rcj�1���$*Q��K��^ZU"��eK,+i��T1!��h(�+�M9¦�X�dw�ȟ/wՈG��4�s���!�΄�?���Ŝ	Kg�ᙬRp�:i�>�Lu�eFw}���`��?[����]�aⲳ�(��j ���.�I���T��V/*:;k荷t!�/�JJ���K�]��`+������
��T�}@泻�W͎k��$�$�7A���U���y(�� �e�%wW�]��CWo�
G��Qܔ���ux�e�* �B:ڧ�S��6�D؅�T.��6,�[��P Z�NSY;_���SJ0��ƿ��'h8笊*�k���C"���|k���sE���ɤ9C��j�!H,� �mF�a�v߅�U�`��3���^�]\#j�f�	M��zy�./�+��=���0�����w?�������?'�!_�.-��o�R[���ѐ���`����)�A��o��r5��0��$c�;_wC�s��v�
f-��)c]���y#n"Ù�������亦�H��?�u�X�?����@g�*u�����s����؛d��E��b���p���v�MИ���E��F���)Ը��El,h�Fc���ʜEi-��}�� �$���8�X3��^��5�̄���_���0�w��r!rGKC!Jd�;�ʅF'_q��%�F\�~�ҹN�U�°����˄��_�k�"HC_���|�Z`�F z]����:!S�J!�9�^i�v��|�+� W�$y�:�?�E��!4*rֹ���A��6菮Ȣk�{���s�󟉵P,Imkg駽I�ɑq �{'*�ï�(��p ���w%}u_�H��$e��%��=(t/F�=��8��N�*2��8���8Ci/@>�!�:�|�@��вs��&-$Ah{I� m�c�K��VV�*�����qj��`[��,���&���0JK����XN�^�Q��T�&��g�t�8�Ł�C�Cb�FO��<=�_�d/ W(�e<�k��r,������^w�g�vТéY�a3jw˂ӯ�f]ܴ0�8R��)M���*��(PЏ�|��^V&Q3dQ��u9�Is�U�"'�^�qi�ɫ�|#8����d��h[l~Y1϶)L��
���G)�G�m�IR��(���Ŝ"v�|~��T֡�7�|n<���{�E�mZ�����9ȁ��-�p����y�Oڜ(�~:����FL��'E`z)�B��?�ƈ.BJ��@�����.#�`U{� f���r���,� �}�n�[�)�ҖHua28�B憌C4�^�O��g�<ϟ��[��*Q�,�p3���0\�MnsWѕ|ւ�=�і?���[f���m$�ȁH��J��2�߱Y���O�x^7,�ς>&I���rD�ad��rw�9"��֖c�=�׿?z㞒,�f�&bb!��"�Q��M���q��G��ݿ��
4&4l��o�l�