��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�v<��m���X#�m�o*�����z5�22�8�G4�x�{[��IW��(X(_<A�&��աW�����T��)΅�A�P���)���0� #7><����r|ES[��~�D $:_R.`
Hաm[��B,�+�*	p�xX��$��e�����?���G��%Zb	 ���5��G��r>��T�CF*�{D�̟�[�$xi��:Ԗ u׳����.x�7���*"�k��c���a�-%}�y(>�hž���4���^�X#�f*g"�g�Uu��7Sh�	� �ƌ��!����盛"��q�#��SN�5>-��=�Vg�M'J�����_;�dH�K!Y�I�.�I^�6^S<QѨP�/t|�z,�廄y�9*��|�`=��p�	���=�~�q�SvH7�v��{'���r	�J��仿�<�w�h�4�����q��K���Pڇ�=ծ�*�5�[��Y��e��@(ȫL�M�ٕ{R�Ϳ�*��ᱥ����X��B�p ���#��uq�/)��jv=��ɶe�Q a5�/`����R��p����~r�g���7 �WH�0S�A8B� 1��26�S1}���� c��^5
qgя��Z�G�]���|򸏤�r�HLx(5nM'�^�Ck���	*��=��ݐ8����@�}�黮&]����U�ȴȍ$���d��&���+�K��*��61�Um�?K�O��l�jA!H�qjfr*!9�k�rޘ�q��X��جGs�ξ�x�0�y7�e�feZش��bT�ѯ������l�#���z$�ʽ-��U>)�eqbO�j��򗙉2x(��"���V�?꣕o�H���Fa���@$fI�8�:�����H���t]=���DP����C#\FU��1��(@�9;��G�!����gʣ�@*%/�^K��:��������ޮS�8�=#�%O@Zay�0I��g��t��ƗF�*���<p�|�p~xjV��셧���JD-,G���M�a��d}S� Ơ���1(?��9��'��7��@q>�{����w�\;`��lx����댠���Aq���>q�dB���JN����.gy]n��C�W��,h� bG�p7y�g�=Y��.:��u��;��\-����!�u���_�fs$�\ �C��!��1H�Ǡ���������>��J28=Ģ�O��;�e���
�L1��C���ҹ�v��fc�}��k��a�xJ�(�5,���"��X_c��J��ZG���Z�	�dg07I+)�f"������1����ۧ���,a���hS�l��X���Ka*}>�5�������@�3j���* #�?8��7���ѐ7�<.:),l��@q�=�#���ZN5��H!���/�~��oaW��¹�؈���[F�V=`�L���R��H'�4H�Xb�'=��Fx��ML�kI��+h:VDT�!n���_[`)_��2�}�.��-��L"��=��f�f��,�h�����,���a��o�	#�{3{x�b�}
4�VI�B�Un��	��[�����{�8�>��	!�qi`�w�!�t�UO,��]���}G�W�����Oii"��|1�}��A
�*ϐ� �?N����L�yX�>�j�^9��sti��d�����o���	�"���b��I�q�j����`Jȍ�"�/���Ż釜����Z���qi8VU#i�c�"�Ԃa6� ��tv�����ɒd����Y������G2�ڄ��	5�@.����X�6�h��*�E'�}��U�����άJ���>@.O��j�z�uۏм����v(���VD�G�6�dd�L_�@��_�(��6QN'<U�#G�`efl�'���Z%�y�P�����?�-�����>��N��J<n�a�p���Oj�nd�n�
�zY��������jf\�b�Re�	������mӜ�l��!����i�rT�;
�P�ES:VNh72+����Y��3�Y��%G:wߺ��Y���� ��]�/ ��㶱�\n���uf78#\���Y�t�V�kjeٙc��!�l��� [U�vDN���o��C�����;	�M���~v����c!4*�������^��C,��К��_вl���w)�V����{1��;nR�o�����ݰ���@�^����[L�bN{��?��fEjk=���`�5���"I4�=���o�m[��������,����<�!�G��2�8�I�V�E����2U�FK�Ɵcń�#�n&cdxDD�t�+P��{�ZK^�­۰��!/g�\{��s�j����Fu�XS��#w�$أ�89O����'N_��0���9�9Փ�Ո�/7��Aڋ�w� ��̸.J�S��o��n
� �*>;��~��=~yʛۿ�K"c\+�����X��|�<�j������P��t��oP�gj�Vn���.=�2eREJ!�ȷpɠD��/1��UkYS�)��B�E�ZM���k���z	+ ;3Hy�8�����R�Sm����0�IY��A�Զv�ӷ��~��Ɓ�T!����\1����Fh��P)�Vp�X�")�9����3h�DuVF��`�I�N�l�� ���S��o���K���FD���6[��`{BΕ"��:a��IU;����9�U��ק5X��8ʼ�0� �m�+Ε4�����\�;��,����z���Cv���HaH��S�B�\�)��j���2�����{���Q��X[�t&5ʨ�t����1#K���+s*i$��U~��4�+'��q�V��oil�v�h�^�4�B��9��C��_�c�	(���:������B�\���2�{c���H=��"�%&���U�<=?26Y�|0���8a�����3�NW�>%� F�-g�����$�]岖H,�~l�'_E�wj�X@\���ω��5�1YS�)�L�?�<�2e>>ްI���X�k�Aqܯ%�r[��0"�*CA�X;��ᄭXMC3Z��p�E��I�sёW:��v�#t��P��5$��@�%I��v.�j��2']K�v����S�Q�Xq	b�)��M7+ZxQ��_���Ǡ*}��]�Ȗ���(-X׾DP�V��?���7L3��q� ˶Qt_�øÚ���[�|e
�e*1������#���2���k�8�|o@I W���R�8�V��X+<N�ȁ�!)>��+�tI`u��OCC��Ʀ�3��-�<j����/�����S��yL�l(p]�U�|v�g����R�_ރ*���C�MWm'W���{�-ꂊ�"�F�z1��9+������z���/��pQ�I\�q��HdU]w�4�m�E��5�.	`���zȆJ��D����Ь���i,Z�{�s�K��f��?��o?wB#,u\!ҩ���X���g�������b��`���?��M3&f�)}�>T��r�\�Q^B�~��F��grc���Ur�*1�������j��	�1����z�;.2����ǻ���$7X���@��ҙ��}J��%t΢�~	�a�غ�9���s������5e�,X?U��)�ƽ+�N��L��x��
H��4�j4��M�x�g1�%���ld}�������d֊�~WB���Hp�!a�ڢ+❞��TP�<���WcHn#��U����*c��k3����� ��q_����˼<Rmv{f�]wY">���;D�4�9���0�C1#��D��z����z�Q���������0�ӝD0UƸ�l㉌�?^Q����gv��{�ѩC&�.rG�)ʔ2�9��Ϧ��V8��f���E<|�S���c��*����k���T/(�G`�p7���_EEuZ!�V�$mv
֣;_��:9�0������>��^�,�G4 D���\�����l;ܗxL2�>1_�Y,�@l9�+GG���pC_H�d0�8�N�<���)����G��Ud}L�ѷq��;}_֡Ux��n��*�#g`�ʶ8[.V>�n�<������e-V��2dT|'�}xZ:w����e��2�F�����3`��3�=��(Q�v��N�%�^�;:{͢��e���Fܥ���0��O%֚Ō|�l�#����6��ћ�t-`�4	ߕ����F*���.������ B �=��O�q$�����hP�D1����n@v���2e�S���z�;��+�N��b:�4j�5p`��"3����Ƅ8j�ℿ�%��)�%:m.�"����ѿ�!1"��{a}�y�˲:!�]�d�T�<:5V��	_B��КQ�<Q�E@H�7Bv���La[��/*a���0o��ل?g�/
ro��:�!AE(#���C,2}g>�ـ�#��n�J��xl�"��ŔsP�"���ZP{ɑɴ�/:��f��y�)3�gaS��B!V]d�~�i8̬���tZ����_�ȗً��g��[G0t�i
�tӖ%��L��m�[S�P|�z6�s�@�a#���V	�,p,�E.� �ç��[�8�ܔ���'o�F������N/O���n6���ê�����Pv]U,P3�wW��=�3j��F7"��:S����#<����ы���V���u�Զ-j�b���a���4�̜��B�k�>P4k)�7؏�a��Q2����{P�-i��%��p����*Sc��X��A|K$�2�#�Q���jw�r�$V~�,�����&ī�S�����#���`:���Zڒ��}����p�c�=��`�	v��J ��u�/�]�")I���MZj:�������m��6eW�eC�yA�D<���?�%���ׂjhOť�NV+��.%�+ýR8w�"_��6"5mBQ	�cU�$��:ۋ�Lr�}i仅�y��3�	�^yQ!��|��<#���m|��ZRP��Z�	�R��o���#��ro����b�qj��n��7�{�@4�1�������֝��N����N��-��d�X���ޒ��N#U�$(��8w}��jK4�yH_$�Vc�Qu΋�Avg�P��N�ܚ�����+yR�[]����G��e�yV��@�������#���o�3�hL�ܯ�hZ����ܽn�@���B��v�3P�hP��f�ͩ�ϺJ>�^*Hź�Z�lJ�ig��U�RL�LY��괱R��s�2�}q���&h>[i�O��X(�Z��kܠ~��i���G��p�ZLv(����,ٳ�۵�7%��@�%ŀ�F�z6\���zO}�@�3��E�q�X�6�M�*�	��p��j'��E��y���F�[F�b�:�����CMKȞ M�d/}�|��VE���ՕN��`�Q�B�?����k2c�.�2��J�A�r16��ƍ4N��Oor� U�>���lߓڡ�nNH�!'�4b�]s�: Mxn�S\k�A�v�]��6m��I�Ƚ)����������6�X1�7lR��i�t�4�����,�>�F��R�%ݞ�Sp=\�L��ة� L��P�{.��f�7��0�Cn���v�Q��@!$���ү��Aڀt?g(Y����>:�G I����V�U� �ۚ�u"���;l:ј�N��W��c�3u:���S�6��6�;T��(���f�T��r���'+�=4�-۷�&1���W��P��+�Oț�q�=�D�/�]�*��lZ�b|/wa b��>�Ci^�x�vЩ��x�8격��.K����a.�<��8%����r~G��n�e�}#JjI�ߛ\R7�랃|�e�� �� �y#�Z4����+�r��'R�@@?�(���� 6�!^z"w��:N߂��?��3�+�A�L�K^P[Z���a���?k������l�"2�NR���b�ʍ��]F�kQݸ�5I�]�q�^}ɠY'>X ��}%d{da��;@�>q~#���RW'��}L^��Y]熀�U|8�ҕ�ß�ǥei[J�;�Gv�?��dA�K7���@�J�P��eӇG�]��8���;���?fG���LW������	�����.&`�	W��}<��%�DmG��P��/�����\u��:�D��*��iK/߂��)F����3���L����&�F!{���O��	/C4+���_�\ٹ��w�OB(	���� d�N��Cʯz(��Х�������z/_������lF��2�an^T��iI�~�G�?VB1T)T1�:8����|��02��xߞ�	mq����f��֨iy�T�1-�9H��ؤ��]��ug��p�������DP;��77���S�K\���v�^���1\��v۽�����sn�Jv��X�S�%fP+WI�����f��*Y��Ԙ�N1)���/i#��l^.�g�wA�@� ��R(?��BLʬك��1l��o� ���y,�9^o��Ek���<Z)*�[9�b2�]�w��S�
��IS�K��	5:��|�ʾ�gx�6�r��%9Lf�]�W� -��Yj�NX���B@o�C�&���f J�M�|i�.G$��I�+f<���b�k�K�N��˘�9�7���>�����ZF����"͛��"���S����ۊ����D;���w�K�5���6G�f��/��qW����Ť��`��������AK�ijI�k�U�ZK#Ų^4@���Z�
���~@�'��������a�_�th�5f�aQ�߅�����xh�eX��=�t�}�l	$6���@��ܞ�����٥�#�ո�,�i��ۨq̷	�n������9R������s,Q�
���2������=c�O��B:���AW��ձ⋒\�����zT����H`�-�8��+H����=(u�ۏ�X��X��맠�#��D�de��#����hh�7rUx�8x7m�ʰ�����$?�,}�	�\�ޕS%2�1Z`x�S��d��4��r���.�{!<��9���b�y"���"'k�
%4o^IN�/���
k�{�o^�6�9n^������<�sX�1SӼ�O��*�A%�u��s��lok��廬��ܚE��PF|y{�H{.�����]h����a��5���������7��꣏/���KV�����~�6E�������Ƚ��P�'�����x�^�m~��Z��,�ES��ҟE<HF���In�Yi}���4ˮ6I���t_�ơ�%c�]��In��!�'Q�O�\��_c�+L</��&��M�����/N�����"-��M}�K��m9�W���@v��t&T�y2\��㶪 �|��kš`Lt��K��7��[�HHW���h��Y�/�ƮX�����`.��;"�eV�UaA=m������T�6t���dC��Ug��=��x��K����ε$�cDo�"����8�9xP~�@6���ߘ��i����K��X��]�E^�0��	�l ��;�]J�i32��y�=��i;����~7���Nz�iT��-n0e!���ߗ.���ƁࡴN�4y=��%�,���k�\��QJ��4�,Cm�Wڬ��2}y�yO�ô�H���:�1hRٚ2�6{đ�◱&�yg�\�D�j�siSl���W��3ώ�;,�.PĎ�������~�9�v�Ե�
}aZ��Ea;,	-\������!\%FwP��B2I5CA�ϐ?�Tn�1�Q�u0��ꢇ�s�<(���/K\=?��(^�赵��D����*�3��o�F����9%��t�غ-Vn���/hkz��k��s�-u���*L��B�V�q�	t��Ce
d[(o/�f�~K�^:P�m�3�y�|�F�s2I��ek���&�[�1� ќ�-��3����͘��01Ҵ�����Dj��U�ՉW��FR��(]�_��)"L�A�o��>�UL��B��]��#���q/>�$"��@�o��+j�0H5q4�kNאf�xˈ�>��]�j��xI���/:+R�ti�򗥚O�]�cp?X�ّU��(݋��XW����/��Se��"�Wp(;M7�*���X�M���Z�K!�b��(7A
�M�m�`��nOa2l�c1'����O�=�
����͞�{ݷ�Qd��%Q~�d7�$�t�j
���d���'������3��Z��sR���=p��S�����]�u� ~�ψ״β���9
~%YB$��48�1�A{���А ��s��)��+�Z�P�ǡFy˞���C���paXlH����iv���z�r�=�̿%�������~��>-(�	Q8}��2j�Ht D(���Y�PL������F*���yZP�̳��ޚQ�� e]r �|9{aܸO���cv&�Fg��a�}b������B^aܢ��GS�J\��	H̘����^�W�~�.�+��!�Eqq& #YT54@)���s��>�\�pT4�0�%\Cx�=خZ�
�@p�-F�^���o��� ~�o��1O#��:�dmNP�d�s經u�Na�2jS���v�l�ra��/�(q� 'V�����
�_oj)�&ٹ� ��[^t��y�-��&�,�\\c\���2c{t�M�|�@�����*��ԇ=6v�x�����f�ӷ���tՈ&Y��7S�"5�yɯl�{�Ѫ���sw/������T^FB�b|3`G�U�(Is��|je��.��'�;~� �m��p��ʽ�:^B4���?�a�&rf�i�6�0�_Z�0�x%�?,ͷ$�����k��D�X���%#J�wq�I|Ή��ɜ6����,���d!0�*ȼ�n��н�&10��5?*��,�N-�O���B|ǒI��mZ0�g��!<�:�ܹJ�ۑRO��_7R�a����ݾ1���;|��oB�)��h�ecمI�d��V�Æ��?�_�H�eDa��Q;�����{��s��7��j>��� h��g
{�ҳD���[`��{�?oi�0}>S�ŋDt�z&Ih��Msr���A̶'�mO�p��Z$�`�c(y�t� c�o����LfƝB<A:QFO��^.h{���_j�/}�HL��JV���w"�9�'8��UrU��8��"�oQN%��$�]��Yy�ff�)t\9�ij0���$K�a��� ��s��X���9i`�	�J��Pq�x-�8�뽕�
���|��;&�D���g��]F��:aC�_��Kߋ:( �L��>��A�oN�ČB�7 O�/^1���Ɖ�(yj>̖#�'#��A�0��p�=���"�m�H:r�b�[b%gm\�4�5W�;��Ǜ*E�]��&5����}<��	e�w����a���+;bbV+�,��#̀��6h�!�us}Y\&�	)�C�%��%9����� �����Zhկnb�O,�{�r�\�Ұ�R�̙��DB1���_�6������K���@_��+��+ULd�E����\Į�����XFԸ������L衄ng ��Co(^�2$i<������L��⌏�,~��\)O5|�6�T��P�_�������ecxy �O|�]vGҗ9�6�)�{���s��he��l!��;m�?a����V��'x�)f���H����No<kro\�ٿ3�[Ϯ�%pD�YIw���ޕ*��\�'�6YY1������%�}7�����n�����u[+@.���gc��v��;�gI�aLqǬ-[��~]ʒ�^n" �.g���-YOuy��Ⱦ!�Pk���r�+�F>��:����\���߼�E�c:�]w��m['6�5�kRMq@ӄ���oK�.x�W2�=�Y�;5��k�" hx�ܬ���P�h���(��/�d��F�	���sc�¨k%�)1�|�f4�C��o�<�p5b�GѶƄ�:+��`CX1Q6�ta5��V�#:=���,T����>y��B�t�Ap>��2R�R�:�7�/X� ~�a������W_�~w^��a�O���9�mg�����l.v��8�������i��)���\<.�H����u��[�F������ǎ�(_m��h��1 ����ui�cY0 lZp��X�%�0��.K���+�^��&\���"���4�Cl��Y�)�>U�����JI���u�7�A> #7bNW6����Ƒ�/�7���~iջG�3��Ԭ�����R9�r:�{&_��E�/�a�c��I�
^$"q��0��e��h����(�5���(#�������vbٲ�Z���PUM���_5W9��;�Ԝ���V��U!��G���S��7����"��x ���Z܌gW��>�+{�yq�d���0U��_�d�7�V;��o@�{�66F�VgL�p���j��?%��4��*�'�����'-�:[��-��w�A�e�h_>թPݚ�3�3��O3cT��.��,fs��
��z��%"z�6�I1H�L�wEh;x�3<-T�_s7�&�٩#��W��l�#������L��`/�i�'��*��BM0 �D�m`~dz�bbP{ƹ��	�5��U��t?Z��FJn6I��V��Z�uZ��пI�Y6����D��.{�LiH���҆��U{V_���&�w���z�z.A�B��{���E"u���b��Q���l9$X)8�j��x��ZMV5|4[�]��g�~ ��Ð�;�E�]��s7�^)f1,��qw�u��[L��Cd�B�HE��\����)��������s������M���F�Ty��O�g:I���`
e�Ľa�\�_�����t��G#֞��oX�Q9^B/x'���y(8UJ �|C��?���M���,V�V�
n�@��E�����Єtok@��l%>W
�nc椵Ѐa��1��f^q7|+��ಏ3[�kbq��9�/�����"
��ࡔ��;�/S���C����?�T�u~9��^|OC�w���
��PS�����bѢQ�(0PD�Xqy4r$�u,�\��lM|�TN��
5�s->��C���`���q��
��´�mR�)�E*:����x��}���XD�ԲGLFF���{̓�����c
e#��.D�Qs��w �Wm����eyI]@ތe�~k����<��0�	bs��ҁ:���Mf�- �=�����ݼb��"���;��ޥ���j�C�1~�E������{ft��2VŅ.����͋#�VI�f�ɡ�\:��6՘�6y���mz���d�'͗����,*$OR��J��O*�����ts}RpNb�@
�V#��;˱V��V-�qcԤtK�v�W���)|���ߋk��.^N*�wp�bTpa@έ�:�-�n^���6'���{�<�ـI6j�$/`X�yG�^C��$y��{�k�U����Uhs�<���.$&{��Q�Z�Ll�T�Q	�Ic����hՌꂇ`����p�<Q�u�GKU��M��؈��	1r������ (U���� 5^��zS�Z^[�+�(�@��ũ<��L#�Y����	���2"+�� �Z�ƒ�ԐrY��E���␮0�l��27P�a��p�-~�bd��N>�J�m.)V�n�-��P�+�A�0W �s�ܢTн�_%pFu��y)-74n(�})C�D%J���TN��5�~䕬��F-���bh�Z(QM)��a'H`[>�e��_H5��a�z<��^]��&cd���a�F 9&�{R-n�1楟T���]���,��y��a�����JJ�ˎ}t���cs���~���t�W��(V�>m��<sd�˔_xM�A{���:��>\�{u��c�Q��B�^>͆2m[W�i�X����pu˘j�����e�����5f9,��NI��l��F��{���� d���,�0n]�|�?�2Ͻ57�f#Y/��?���+�k�JM-� $���*([��Mvפ$������i(w��@Y}���XӰ0���$�tNHt�ҝ�kt�y\��Vq����/��P�]i9���&�Dv�⾨i���$��X8ȸ����i���jq�<���$K4����M�w>#�Z*�z��v�-|�BM��)#�Ex���n�@�U�����(FQH�ٳZ�o<�#�h����oخ�{*�H���yu����F%�-��*��G��+�:��d~D�D꣟#�F։����![k��e��C���X48h���+�p�#j�u�����T� d�g%E�J�u��	M�~FZL�f�3�!��J[�W�������_Qʸ���QF�m�r)9��Wߞ@V�7/�9G�r��L��oC̕Ju�V�w�V��Y�qI��]2���CM��L��&���Y��2���A~N�^�IdR���c�Jq��Kl{R�&�'˶j@	G�zD�Iԇ .o���qk��=�h��������D����)�����k�jԼ�M��G��z�fقZ�@��&K���&(Dܳ�c�vB��j��
9�$�^F�w���W��H���-F�n�2[1�9%���㯮ޞ���6�����H�QC|��VR-%����}�pV���gt�Z�x8��#�� ���T��Jn��y���EfZ�M@t�����(��-@��i�xYbw2lw�[�5�7���]�S��� ��V�8�2��2tBG�����]h�3���/kЎ,��^.ᐪ8��F��k��:j�B�\�]1�%BAB���Ip���hWvP�T�Tsu�fs���Yu��x�	�ݜ�
�-��T=N�o��:j���Rkl������鵰Р�̝N!d$�\�.�����,��y��Šh�sȾփ�}�Y��%4㵮3���3b�t|l����w��v�δ���d՟EiLA��˥b߈� �a&^�`3Љ�y�=�|�]���YO��n��i��5dR��=q��h������hW\g�����W*OU�բS��:�=��R>z����X$�L�������y��O
\&A�!>�\��^��W�Li�9i��*�̟���(��	�����=l�eo��^�!� ?H@��&"M%(�\�1{�xuN`LBН	�U�c�;΀[ݡ��� ?���{1/~W�o#R���Xn��c ���
� ܪ*&��j�R�>I�o���	�',>`������W��ٵ����rJ����+���i'c���ӱ �#���#a*y�����[�Q��A�8a��K�N����9��7ey��Ć{Sұ&֟-1 �D?5�m���6�!�t��l�Uh�l�ﲶQvL�,�ɸ�h�����K�.�zA���B�*�<�����,��>iA��b{%i�߬��f���I�ذ��`�C5�(	q-:O~NZh*$ź��m2߃���� 1�Z�1�+���!z�6h�0�mܠ@M)�1K�s2��f�E=غY�%̌*��cn��yjbrN7 ��Mj���	���Pkp����y:Ҷ��x����R�s����{�.�"���� ��!,E������,\#ը���p�����46��IU~vO��&["�Ac�?)~�;�]�C����L-/N:�c�k����;�w%�5=��G�8&Z���Q�9(K-2Bԛ��0H�H����Qd���Ԗe5�����=c���m��7�l���銪D�p�|^@����X"3�V�5:�!�$>��>�����.�<�@�~� /�����?�$f���*�%MLɨ;�A��#!�qRߒ�	�#V��y����+8���*��a\���/��n��R?ͤ� �M�S0A�m{ME]V<'�o�H<�\�K�K�b8(��A���(�{C�� ��K�W�_[����y�A�&��Q���~�,�$���AH�j{gM�����w�'����W#���:���q�+t+�21ew�*�Ϝ�8�'z.=���7'��DO&$������1��f�,��4����l)�$�]q!��Z(M�t��� ��:0���역��y�ke�Dwv�)x�zfD�|?Q�Jd	�5�����31��bv�QO��C�"9����OY����N��PwP�T���v�"�=q�c��*;BØ�����."��Ů�i�K�8 �m�Оp�Twg1��.���}�\Q�GZ%��M{�3��7g��1v��n+�`]Ӆ6Q��v����wH`i��i!�	�13U1@LWxzm[�4df+c��N8���)k��f�t�ve�f���m��<�)�����
y=Jr4�"����K�L��K�B��78|��	�x��|�5%X�^^t��QH�e���\Os��_{���g�N�c,lO�j@�$/���#�6���"����|�)um����H�&�W"����5�\�ltJ�K�`k��z^"o�j�߄��s���W�e���UK������^���Xk2�x�^���T�Y/+�o�m�Ȭ�w�n����Z.��{�UDW�m�D�9d�H��w?MMj�")�xT�kW�y�D��%��C-�=ʢ�'��IZ?@Tt�W�w`.c�{SO�����@C�b��l��|��`ͱl4�n�LŽ_Qp��a�,�����d��r��������w�Q��f���\V��'����8�
�'+ʣy���{��^��R�O�7�'ujJ``v�
�>�J8�d[�z����*p�(��1&HK�;qa�1��M�)IL��n#�k4b��I�y��w��Ĳ�SթT�;�3�i�N	���w���s�:S���4��g�lG�ՇŲ�N�u��\����,Ņ�S.��������7UJ�� ۫�`� ���p�8����ГQ�Q��l22H]ͷ����R ��W7*>��Z3��J()ړ��~���mSL��R�y'�ԛdq�a����#�� �T�AJ��9?����Z�V�'+��G5��h<&���nr�����PM�=eݒ�bSy�ʵXhQ���9[����eʱUȭ��Ӻ|9k�����25��;�Y��U�E�i&a�8P��X��]"���Ɩi��^��Imd�4u��a|m���8e���&}���k���"�WX����G����#��J"��-�)ס���~���;�O!��J��X@_���⽛��jx�Z�xO:��l�A��)�qP����
 #;�q����u6E�Oaa�c?�s��p^_,�EJ�;��8�tSU��������@uU����@�`�9��KR
Zm9ui[�G͂�TVw
�I�܄|'6x�CۿQ�zF5����Y�� ?�Sķ�@z;o,h�]>�)�ch�Y�Sŋ%bbֵ�j�i�+���@����1/��kQ���+��tuE�����t2T�Q6h��x�g1v'�Q�,x�t�������[���`��p�g�hV�F�H�V7	F��މ=.��C�0V=
�߷����Џ9)��e
��n�ι�3}oi�����9]�d^o�&VV�*��1��)(�@{�'�*}-H�h��=}�Z�N/���@|�w�˸3�ԝ�Q�x_Q{X�c�S�=�#�#��`Ǔ���T6������j��"�-�?;S��$�I��
�g��@A�~<�O.���bL�`�ZR���{ ��#��ߥ1�i����}ߒ� yayŰ�#*�e���J��ww��JP��{��.�oUV���Ͷ�V2٥x`D`Ԑ۲�5�,}1���Rh1D�q҃@���Ȭ`xn]�Y��.4�u<e�,�sz޴x�^�)Z��;�>{��ջy��;M�tOD"3X��z���;窴0�A(�Ҷ�4ލ��a�-$���HAOk{:�4����G~䨸��l�����S�����n��%q�9&�rK޸�-7����n�vJ��m%��]��o�RPz33C^��C��i��ѱ����� ��r��H7lq��8�dRE鱯�uI�oC�F�;�c}q��B1 �$)�������ωJ�Ny}3����,�u��d���1�1������G��v�c5Z� ����VM@��J��-@�� �!H˼�V&�;�#��r��KY0,,�\���JEY̐�>Ң�iZ���$�(:[�DY\���;�~c�_j��\�>[gA�q����k1g�t��e�X��~��I�����YY�����V��1̬e���1#���M	�s`�\]�8Si+�;>w|�9��w�d2@p3�n����>Κ\wa�]��G��Nt�0C�-�G�ݕ�K!�b�͋�*V0��\O{v�(��'�!Fө�>�\�y�|&`�
�K�e�W2��Q��1�cQ�p�vT�� r|H���lU>[d0�89J�)�/z,A)���+(oa7h#�A�]�O��[�7�������c}O]
Q�{a�mE~�4u����(5���Ms�(E�9O%މ>�ET7�'V��T?���p���!��'L���"��s@.=�ע��	�qi��.b㪾d��A�V/@��r�X�H!*���˭��	D`��ϥ�����ܯY��20@�ax>�m�}9Ƣ�w3V�3�K���'��o�E�ao,�hL���C;��/����U�,�Eow��,�L�+oh��r?֋k�Y�Q;���@o#L�Z;��]�w���z��4�y���^E�Q����������%rMݔ�:澙�~�Q)�7X�\��hB�zG��j���)�"yz
�s�]Y��k>��ۼ��K�7�2N�x�u0V�~�(`�C���[88%f:���p�L�����I`��A��1O��:	�]��Ŀ����1�	�B��g�tg�7��"ҿ�^��j��H��8"�M?cId��Ī�E`/�~�b�1�o��;>��e�o[���ޔ��f[:)�Rʵ�!y�Gm�\��o҅H)�}�ϩ�jU�Dk
]��/���a/��}��U`���ܬ�#=�xY8�>q�C���U�\����A��nс�2f5���g��b�!�F���gHt�NN��┥��8,v�֒ߤIקƑ��I��H\ ^�%Y�Ҫ�j�p�U2�쥍p�y�,t�A��5�Xȕ�.q%	"\f�`}!-�n��f�@���NɣiHA����p�|���K{]��`Z�.��s���"����n�%�W|��i9ʾ%�Л�����=���8��x��z.�4g�Z�`�0������Ώ^��~U�*��ZϘ�����,_����xH���HI��a��\�/�j�Ԓez�!r�$���!�x=Ζ�96pC#_u��b�\h��e)X��6x25�:��*?C���[��l�3<�(6�A�붷"nbܰQ����Fޯ#����e�N0�]çA�7�(sa��}8����IK��ߔ���}��(�.tr�zd�����0�T;3Sfnb&g&<+��~�J'RE���qҿ�J�p�s���%���))0 �\��8Q��2r���#w�ӌ��c��"��r�Y�Y�y]ߥ	/��|��q֑\k
�g�l�P��ZTh;{��~~[�s�Dŗ2 &�\Vʊ�}׻�~�n�l'����#|'^8�h_��
�&��;:��w��c�J�����0s�'�����p����DFv���<k�����nہ_��X��J����(ݹm[�Sp+J��]p.�����нd$;�ي����d��ێ����3�u܏��w��@�A�.?)�qݥ��3o���^	=���J�����x�@V�*23q0��� 7z�AQg%�bF�O�P-�.F�'���6i^���{��_!�۞��9�G���Դ����KW�%� a�uqy_�%�"��ݺ�
�A�YW�<�d�k3�#ͯ#[��%�p�'�$>pm��S�K�Tq�wfm�
e3;�v��_i�]T��_T�[��6˥>���ф�qŅ������!Yl��pc���:M8��d
�9m��TQZ���6}_�� 0�c`x��YO	�qIv��Z��䟗��"����=	4�z������F��N2.-��T��6i�,����Z�d`nw��QP�c�N��A���{J�r�Ы]�)�e��'��5��MG�	'�;���Q!_�Nu�Dv.S��P4FJ�~�7���:��h��mY[rp���j;T����J���~B����BX���!iGa��d�ѭ��P�C¶<�jًd~�dlg�k�W^b�-��Ӣv@��� !���^�k-�u\����+�/��]�/�F�I�M�	�3.�.`?�6:��Ԕ� ��s �bV�h��t�\����mRz�D�������������TA�m�N�hUp��9���7��0���h��M����)����BeU�G���%����#n��������,��m7�U	K\�SA��V{��	�s8�*9�^�}�!�:�K��D8Aq+>΢��q|�z8�s�S��Xs�՚�g��].�)]=��)�A��V�ݶɊ�e��ڲL. �A��viO���~����8)y�������lcX�k�FG/>��8��r�������7�v�*Y6[�hi�h�5�*7�C�i�O2��<���7�����cO3D|5DHJ�JEbX��p�$���Tq�����\	�����5#̮�G0,�v��v�z�9Q|�_��K'[`�*u�嗫_+7�RK�=��s����h�T�����3al�t�b����F">h�Sm��fs�QUPEQw��4���?_R+�c)$�5.x`i���
�#���^�z~�Z�2�(���L�=����GJ2�}4_����_)�h����s������N��F��W���+vԤg�A�.+�+�;���Vߥ@Ӓ4�x����&�Z%�Àđ�{����21�	�&��E�_��ҁ�㚯%�0�c��s�⍑�X�SN;p�sJ7������Q养�eA�,]ց�f�~/�j��eS�X
�P> ��DB��b\�䏝������xpf����Z�b��e��1��]	���~����;d>�W�}��Eo3�9��lTz��$�% Q���S���p\�;5��l���'��U�Pkj�� x�<�I�K9ʤ6bȪ}��$�g.��ʙ�e��g�C�_V���kt4 �5�7#\I�imG�"Qf[֨3���(�1�E�0^��#�|�k1q���/0d鉼ׅ�Ƀ�@�q�!����5�ΫgqEiX:�"܎�GW���1!X0ΐ���siih8!Z��yP�RUDc��y$ϩq5��Ed/��4s=��g�8iz�ם�u`����5�0֋y���$�q�X?���TzUx;t�h����n-+�T��~����O)5$ ��t"S��6D§��Z�$��4�S�z&����
=}��13��:v^�����	���}���i~���4>�����Zf=�f#4*�
��SIaKw�ٴTh��`?��p@��	�u�� K]�9Wo�) lP��'RG6t|Bߌ�KB�޶���80,2�6ۘ4��un�<?�5����T��ҏ� �,����KK�;�%��J��4�
�<'#����b8e}�00ncc�lB@f�J2s5�5��eb W�K����K��>a����Y�W�"fҋc?ņ�7����XUnp�I��=T��4R�l�{D�eA�+h�
^O_/�`	9��a�J6t��;J&O�q����A�j��lP±�c�3��k�bz. 7�����3�4h���f�Ϛy�7�ȉ���7���e�g�d��
���.�\'i���u\#��1'�b!0`���T)gt��C�^���,���M��O���;�_ �>��Z��|�?(o�1��C:�g�P��Q����O"� VL5���e1��#����������}#��XݐΤ��H��2}�;�,�r,W&%<�:Xגmn�,��W�S$ ,H�JK�d4_������/p�G~;��H�B[҉ª��"���:[�Xh7*�cR7`,[P���r����28La�q��AŐ/�����4*�dy*O��P|���hU/;#�y�̧�Y��ROu���?/3V/ԎEd<�+�.�N4]e�~���A�=ԺKL�s�sa>m�t��&b�څ�@[v ���HZ~�����]�)�b.�b��Dt�n=��޻�����oȆ�5��Y�T���Sf�g����\i0��q�`�t��]�[$� ��[#K�
���'��$�ک)�O)?�4E��[�d�D�Ƙ�gXВ�!g�g�"V��Ip��x֪�`)02�\\zYG��lx$E퓔�~0�8�����v�u��"Q�㐮�^MM5I>q��^��d�Ub�2ev�j}��b�lO�Qle"���Dh�e�ČѥףE�wb�9q��'��X.�U��pؤ��
`�H	P���H�6�@g��e^!���s��#���q\QU�$�]��XS5�	|��6�T_� ��2�͞�/w��f��8�%ZCe�N�?�R�ˡQ~�q�a|
����0E�l_���rNShl,y�0C�Xi<'S�3W�j7����Eaz�CK������Os^#'���K9��良ѣ�j�?�vC��";]fg.�f��	dFn�s��5	U�b���>3�oT-w_��x:�7v$,����)D*ǆ�FڸR�/:^���j)+j/�r����dP�>ۑ�V�$���Nm����n,��ِ|�V❀ ҥ�9�6L��q��̺�G��{bR^3�]?x�>Z��Ӭ��������L҆��>	T�
aM��#���;�O:�O� ,�d��0����⳷*,L��\Rt�k�����TC�b��s�&�4��?}�Xm���D�k]�H�_D׵�^q?�PN#��ȗ)�0GsU�F4L��9!�q��9\���n�����sHο�t66�'�Ŏf�	�(��(U/H*��`��g����7G���R�wo$������J��Z��,�pa��4)+�ɏS!�y^����ŜE (jJ{���j/>Z|s$i�Ց@ �Q�Y���tE�&ǵ)!�1�md�ڲE�N�CR|���O�;Q�����_�����Bm�~mZ^{JK�bAn��͢��m�t-���G2��k�
��6w~<���<c��fRRN�T�Q:�9Vz��g��d^"7�F.�C�{�Sg�%y�.��O~;P��|�LD�;W��[Up�*g3߭=�Bb'�{�o_������#{{�;��u܆/!�۹{�ۤ��V��O�\�D�z�Ӎ7ž<����^0�ea;Ѓ[�}�oT�d�=�"T��Kh���A�d)凛ڀ�WM^J/b�2inF���]+2���/]�2����k󭶫AѮ��h�-�|24łq���|~��Uֳ��do`�u��B����p�:�פ���Dk�]��g���J��']W �����:|�� D�ń�����!��7x��6�BY�8T�#��3��u����5"�t�;xp�m���W`��p���|l��mr�0��
�A�T�˾=�}���
ٌ2��� ��k|����x��4n/)1���q��lJM�Nj��`R�U��l7�Mˎ ��G�����(n�FsR� /Q���ǹ�G���j΄>�e��]W(ź{��z��Yb��z!�Ǚ;�;�B��Ǭ��؊��o,�碀�CI�������~{u.�@|ac��T?Kj?�k_/�|���)����[����6K�y�:��!�ɬ��A�Ő�;�n��e�}�+�d�����x��R�쭚�W=��N���\��KJ�r<�U<?�G�L��WS��)���"F_�Öm�v�Q�+<ҙ�F�o4x��+k���U7A�m����=��*
�Kpr��t1��T"	� oؗ�WO�D���BH���h��.$��Z��W٬�����j�d��X������6��ܔ�U�#�(x-�ƹ�>5�"*�d&D�Wj:J/@5��|�W� �"���}cab ��O��cdx��cM�X�q*c�Z*2ڗ�`����B�t4mĈ��v�f��8,��!�w���������&����K2Խ_�9Y$�E��o-���G/zIOD��z��I�����duc���[`��;EA��Ç�"/�6 �G���8�PY������׳]9T���Qx��Pi�<&�{�����~	���l���x�e�u�Ib�$�W��|.�3\V¬��t��(�u���O�]����|2��mc�7F6�^ClȨ��x5�[���U�P;JYy(�@�8�S��$\P��BZ�F�&��ޔw�P���Sv���Rȏ�u�� .��������̥�XJx�_��t�=硘��.{�Í�ۻU�&#ۥLU�nƚ�)+4�:L1C�_ׄZ��Lk��W!?�_1Fp�.��9�DB���؅��� ��v�nVҸ��
8��C�D~�D�	�,�T��D�M=��Ă(�R�0�	���:q.��$M�������9�(Q����>��s��r���۱��I�P+,�~[�#Uz�)�o%����>I��X'���OǑrxb�i�Êax�9RY��.���Ǽ��n�%&K\��1i��/�T,�tkO�G�}M\�8���I���#f����[w��r�6��p�e�.9�zn;�p���9!Ҷ�
���]�c��.W����M�h�B�W��D�IK�.�Tu���/�>��<I�?����?��������O���Ԟ����)�=��\ᡯH���O*�g�/4I��5�vLF:���r��q$#B��Y`����SV�Q��������o7(]��y�5�׆Z��`�7'���䪣�J��hc�1۷f�B��=�C�Z��	%�^,C�{3##(\\W�7̈���3TB�r�~0:�G��),��/٢�1�4�w���=0F$[�A��d,��)yO���
1�9� �����bX��|;�Q��ߊ�-����%�ܑ���	�Sj-ܢn�Qo�B�l?)k�ݩS}��K��C�J���\Obc�P�d��f��jFҧuC?��l��R޽�wMR�V�K*�?�[f$�9I�^��隧���o���G��YR���p�CW����#Ӧ/����|��K�X� ��A�!�gR^_�p�FT�!� �kvT>�w�L�?��l<�k�oFeU�A�hV7;���H�����rW��@�|����N[de`r�����8�e��]�+��^ƖQ�N*�Z��v$���%_��d�K�æFYU9XSs(����B��̤�������tYm�žr.���	�a�"��	>$�J�8O.a�u"��zVy8�s�_N	m;h�E��X>G�h�2�r�8=�@����P�Jk^E&�<���� ��r��<�ix⣗f�z9vںDLr�UX�ԭ�O�5� ������}\�Or�r�͑�PH�N��	�;z��x��,��N'���sEZi�������G��n=�g�P�D9Qea�ʉ�f�רbv��}�|�r���1��(�^x#��
��t,A#R @3��-�7;�&��e�/��c\_���(:���"�m4� ��n��Rq��f!� �1�5�����ZD��{\�}4ݛ-ү�c{k�"� >��I����#�Gm���N��'��7�
j��HJ~m���{a}f�;���l������5c$XL[��Şt�js�,�r8�{��~����3�gߥ�5KeG|.8�	���=doY�	���6�Ǎ
��_u@�Jxz=Z�G^	����9t(���ފ'��]c��>���w���l�2_�wse��8�6/=x�����1򛏳V�� �x�6P�Ã�l���K�&���wr��GΏ��^:�1ї��Ih��|6�C��C���(��j�\u��h�`8pȯ��d�A�Q-��5�e��E�}���a��vr��'����Aj�7h�Mj0`u�^|Ç.�׹��2��x,
y����ҎB���ա����uh>�@��B�f����jhU����M�^튀�$?S�5�&�����׋�������㾱CV6E�[�^����p)]#[\֔f>��*w8n?�(q� �1Y�i䙉��d�sc�Kq��ܚק�9Nڰ��(���kJ�px4W���;�qa-p�B���!��X�!\�bZ��f��/�儃���޻!6��:�S��L�P�b�}�%�U�T)G��E���M����W�G(�_�H �q��=J@
����'��12Х��taD�՝x�����S��r��)��4<u��L�}�Wh��V���� �='�L�V5OQ1�CtG�t4��D��䏥N� G�X�PU��cq�s��������~N�K��6tB��0dv3*��!-��p�vŻ���n�@�X�;v7�'-�H�k�������i��Y�3��t#�,%����$%��Id43�=E��4`��|���#93��!�>��W�aIO/�����`%&h�T$�B~7<�
g^�F���ڸ 1*Yf�)�RϳE.'�Y�T��{G��ס8��'��џ��`C0%���f��M@�@⇿n�����@w������ O�=_^��;��v�$q�8�{6D ���vZ�E3�j��m��hW|J;[?&c:�{(g�"�{��aiP������d����Ebb�2d-���Dt��o� '�3䣣�&����RX��qv���2aՋ�W�?IP���r�9�(猺KjҲU�!��qBiD�R����1��((g�y%6T^���\G�ۘ�����b�2�k�rL0�$S�^"3��{�;���UF#Yx��tjRE
��<��{�#$$9>�����Ǚ&���A\����<6�q]�+�K ��6i��X�kw�j�c���z��!���ұ��
7���m�r�����.�'y]��1Z�XWq����^���T���H��h	�Z��6 �8(��5Ir5SYD��t����~�l������@x�0?)���4�P��,�:��`�q�?�Ui,���)�N�w5_��S2�ng�U�JL���ہh��<c���~�0Sś��ޗ�x�;�УdQ��H��z���t��mJ4��E��C�s�)�
$I2����3v�@,�ji�3����T�/ԭ2\0���T���(���ՋpF�p�{vW_����c��׽d&�`'���Owv]y�=������iEsk�c!��� ;�L������.7�PKJY����N�}�p�� �o+�2Z���[��r�T�~��'Wɳ���w"b��鳮K�m�dho�>!�\É�oC����au��M]G�މ�MF�N�6�9`��M"u��mC77�3�k?���v��P���#F����ع��`�Y��_
p�=ӈ���
�y&2"���]���rJ��X�T�,c�(+i�&����|��m��Q�nv8V!�������c���O��v�x�}z������yk�J��I�'�����c_腗Ier���E�{����~���6z��I�epv�1:X��Oɬ�J�(��D�u�(l{�Ť��ۗՆ���싌Sc��p�$�)v˒V���,4��e���6P�$ٶ�˧�E�X� �@8sZY��)���̖��^�#�jS�ڃ𴾟��\�<�r	BoF�-G�ُ��]�1���В�2X�ui:�׆��)�]�䄯���H��=b���̓͟�GY7����B(�Z&Q��t��}��i����]�?���(_&���q��?���Ve�H/N�,��~v��(
��wR\K�~�_F�}P(v��b�j��q���00�#/���ЗЀ[�sȺGu5��|5%�&�>l���z�����A\)PX��I}ӟa�t�����i٤�G�5q�s���
ʫ�!��<��I�GL��&��c�*��
d�ޡ�ǵϋv��W���]�����}�G���,�w'��/���������,b���An|��뉫��=�V�zȕ���o@�������&|v.w7��g�����Fӎl~ǃ�Ō�9:9&&9�����b��u��:Z�E��/�,4��D��̔�E�3�Z��JY�Y�x:|�*&C���vɸ��_7&|g�I�|U;ʀ�!�-�_�8DH�������y�y����Ĥ��ttn��am�x��[}}@1�X������%�\���������I����/�pA�٤���-�suL��W��[�RJ����WtI�&�wn��Tڬ�Z��k"Z7�K�SoH�Jarl�A���4k��?�&|H�H�p�v:0��6�W��C@kꈊqj7�5��'�F�I�`߿:��Ue�@�>Nb�>����I�������D�c���X2��ȚX����� 2�:[��5+��зbd���0���^��-٢t�P��;��1�M�����,��_�~�Њú���!:�uU���gV�5M�+�����{�zG?q�I@w�F��$�am������x�6@�t�ϭ�>�9�>1��%��qI#��n�-��U����ԠO�B0T*F�'���㕐��a�R��Q��h`�T���55%\������4�::ْ���P���n�ky�'�@:�2d%u+я�/��Ac��IMSqO�/
�ߔ�����;�BgO�s�)��oo��2��p�j(��E�9�ϢM;�6�#64�W���Ij'���&z�,��f%��K��?���P�M��q�|oǸ@¾�.�1Ӽ��uhm�uw���xu����م�JN�����>����v7-�2���d�9�!�p�!n�_��RAo�5���WL�ؿ�sw��#8sc٨���&�\��,^��4�-#px�QZ��7O<j���Xv�M}7.�m4-t����O�6e�&�qY�N��`#G2���eq�>�8�0�lv�)�a��h�?Q�v���4t�����"Bv����Mk�3�>�}7�+	w0i�E��)��G���I��[�nb���Et]V���[S]4�|5�*f"Y�_Ʌ���pJn@H�&,��~���<��zHvz�o��֭�`��pK}���1L��/4*�e�d답��%�|8$k����f|��´���gL����YQ#�;�Lʦ�d<��&�g#��6I0�j��|ol���1�=��P_z1�m*�Ԅ��;9��{��dU������"�jВ�a�*��(:oI��L9�aX�N��o_VTq:��$����F�P�(�ژ�'X�;�xz��kD����r��mr 6�n���/gs�,���J�v\�����*�Є��b=�9J��t����~�?�9���oCv�p���*+�����6؝�R����W:QC�.���~$�kFCy]H��*��կ9K��+0y��!Ft��O9��s��60�	��\[��dU]��4�-�;��d �,,Im���1��v�j0;V�J-]t����jz�oZ(H��@
<���E�YC��dz$g�����Yq������?���-e�y��y�O?dG!�LC�RY�� 4�s!�E�`ndySK�)N���x�L�Cv��]�j���R��@��&$�4�� ����j����R�y�Jqŕ��J�AsNzQo�Ƈ�4���O�$c�3<˧��i�O֗��1��� �oZm�P5��OjU)G.�^�5�֏K��+}nӒkD)yնS;dw��9ͺ�����������(���}�v���﹃��g�J��80&ܓ�&��<jz���k��o?{���z�+�	2�[!�����iټ�v���O��H$y�����c��w�D�*�����ErZ�hR�Ev��7O�� 	n��>N;�,�\e��G|�j܆�D�D�t��J7J�����te��P׸Z.�P������0�C#�4�8�@OP���6�q]���|�c���SӖ���8�Gm&�g#��9�&�l-��q`�fku+{,0r������9IX��R���,2k�~�Q�x�Ј)�sPɉ��W�p����?W��BK�#�Svكs�r&�.C��x]�r�F��ӄ�i���˙g�/
�1ˤ�fsi�t|F���oFl�L��r����HI����ٝ�J`�9��A�+p/2v�N.~2�~��K�|�<*@K�X p.���s��^�CIi�>>���US����"��N(�H^�1����њR��h#�'�̴���W� 5�d��5���@�O~�j���9?L0����0HS>�����)�(� ����\�ɅR`V��b�?����{�&��i��<�y$.O�Zt�O��' Y֤phη���?ݤ25+�[��;i%wru����F�ЩxˀF�$���G��&/x�
ݢniA��4��$��w%E�`K�( ��hM�^	꜌h����>���_���{��V�[^t����iDG��_\���`&jF���<#�_�DŬ>И�R��^� ]Q |��.�Co6��-\b�)z95��h>R�`�W���(���DxHB�{�%>���,G�ze��Z�/��c�A|s(�~�þ��$���!~����	�b^%��b�E���C�=�����6EF�[α�h,����*�މ�l�����e��8τ�܎��Xuҽ	��p�T�]��"�E��X�����b�� 3Dޚ�#�:�z�'�[0	�����+��H5ʴ[U�Y�I��rts�y�?�vc�P'�k�ƥz#J-5���R"��|2������k�"�_�������P_�쒔��������"��p5D�T��'��W@3a�l	���VZ��Z��r��J��1�l���de6^T	���L~���I>]�ǜ��ܠ�tL�L���VSW(+#�$��
�ӄh��x���O�DƠͨe���} �war�on���|��>a���i��fʲfW:�[�=�:yK<U���u_��>�	K:Y��:ԣ�z�I��N�	�(af>�q�}�0��f�:�f�4��D���@uc*v�$����4P����e��������g�z��n�9P��w��x�|����?y�-��m�hc�˅!�����R���'e�v��(���{���b��1�~vpk���a����9�P�p*��B�V��A������M��t@:h��s����ŗ��'J�����Co�Uy����|Y�
b�����9�^K#���ԍ�� Dؠ�TW�}��FrnW�rc��Ա8%L�NL|��X�Qގ��Kp�G0���t�RA�bp��e��AJ�6sv��3���
���U�u�W��҆�R�dF���h��+ϥ�����cՈ"@W��(#Pw���+pޫD�����T���oL�>17j�Q5�rД@l���#�[�X=;C���):����,�2��y���8jŕ��|3s�y�|M��hLs+���
�@�]N�O�S�RG�H���%gIܣ�fͲ�D�N������	����V!U�E#LD�.��l��I w����0A����CF+�H�Bal�.:2ͼB��ݓ�l��X�-L@��S�~����_�xՔ9vI�L��<�����E�4��Paj�3��HL�h)M���nI1㽝a*�ǬTB:_8�vط3ΏU��Y~k�>��bEf�E��!�85�{��H�����P@mA���q).�,���#`.�0��9n	�.4��X�mQ��fLh''!l�s����_��Fb"�aܝr��å.�̪h�c������H��u�p��G�hk�<a�5�˒�?4�J�=�;�'���`��N\�g�Y�Y��5����f���E&�W5�U�EO��g$_m[PW�M1k���2H4"N��7��=|��m��P�����hq�G�4��������C��l��^x�����&����,9h+��	9�i��[�c����Gl��Sǚr�J�d��AB\���T��4l�~sƂ=���9A,
HzJ��{��9V��Z�(�y�ohAe:���N�0i���s������o��ph��,�����h�D�k��]�R�t�¹aDs�y�57��o���7�A��~�4��ʼ����%�y��� �Ŵ^=bO�L� ;��&?������	.`ܣp����5�ö`YB7�"v^I��\���w��&ȿ:�u&I������{`�C�q���:��A�煞��j?Ъ=L*�'H������Կ��p���;M:"E�\��O	4s|N�Ψ�����@",\��+� ��j���U+³�L���8:t�h����T�����2�RQ�i˦�@���pi@��(W�"�2�x�@����L��sKeU(5�N((#AU��,Lf�4Qk|QF,ָ��D ����¶�~R�O���:�Ft��7�N@��;��ɵ��IF9��V%�1)g��V�}
�K�#�vN����t	��-�+z.d�6�%��U��T�p��?����؏/��)sW$������s���������k9�e;���@(�_�,�p��zT/�u�]B%]S�H`q/��
8�2z�0�]L3�\����2�¸�d�6M�t0j�Ә���ߛ6�ݠ���x�p볣Uv��|�Q	�uӝ�l"i!�Bw���]y�B���&a����Q\O]8 �$�"1��t��ӂ[s'r����i����-�8h�J��ĕ����SV���k��-BC���ae�%E�����)<�(��J��m 9�J�N7�$'�5��q)�[9K	m �hf��6�'Z�M��b�w�lV0�����#Y �>�H�j/8/"��ߌ�B:g6Ă�H��ۤ�Ȯ-�w䍓�V��|�+׌�h��{(���5`��������,��;����<)��3d�7��������g����G��1o��HKƴ�*�n^��ѽ��9Vv	r2���[�c\Q1:�Q�/��(:t�I|quV7$oW�΅^�{[�?��QN5��->A`�l����]�uΔ!�h��Ƽc�)��8��\������mS�����cd���zgI�b3�+ !���HH��z�?�D1p���M���Y�m��'�V?�*�q|oJ=͎Z��K�Κ�������S�q�L6])�6����Pu~W�m�����T�li��]A���(�R�m[��o����Gɟ=����1	_;����Eu�&�$*&��{$����|?F鬭�x��T�C*8=$��ܠ��e�ף� ��>��lq��A����ȧ�xv]P�����}տ;ay9���9M��ֹ���3�S(*��|��E5d�S����,O�{���s?�Fr;�����(KzșE��%�/
�;����)�e��a;mǀ�B�A�x�=P�J�x���hb�9�Q�=^��!b���#O�M�.�D�tω�n��zeX����6 �1�x��}����:WeNq�38%�^׬�;�5f��5�o� �Z�Q�.ێd���A�H´}u.5�C�<�Y��4�!�O��a1�4��.87�_�=��O'3+Q��rG�i{���G��5�a�zUak�p"	|�s �����[�Qd�m�^�@ܓ�b��f8�4K���5Z�7��J����u\�*��8+3��1w�ʉ�,����$��N���5H�y}U��ΌN3��)���FVщV$���P,t#���/�˗'e_UX����s�ω�gg�2�C� aY�FJnG����� J�h��.挅ϯ�,�~�ȟ�8�N䧈�*�܌-�K�,��ש��0��e��Pρ��I����9}Ku�d5���]rME@�����KD�L�!͋�t3at)M�v�U�>5���",ep��^����`Uy9�X^��	��!���=rJ�/?@�TX�O���6[�5)�AᔴH��MH(�AEs����WN�>A�#���x���L�	V@�YM%������<�i*�,<7����`���lnCMӿ?)Hag"�[+L?�_w�P6#:�f���X�/o��2��:[�q��^hx�h^���-����1U�T�bDA"�*��3'�ؚ}�T�PA�J(sWaq� ���dr���]%���P����#_!�eXBc�����!$�I���S}҄�ݸ�Kѥ}v�ڲ͛��csP�|�X��%���we�����฼/���b�k�&�_dq�RC)}]�}�X�0_�*1��^W�]����5_�!�`��?��+�6{����5Ł�W���qO�]��!�>(�:��0���'��$�#K UUt�8USs��.�\��#����ki��g*A�Bڕ��nS�!��椥wm#$\��L�W|�lJ����7�[����'��q��������y���j[P!X�k�*�������#Ν@b}���c�C�ؓ��o���Js��QG7��{�K��_�䧵�_�fd����F)J<>/�
�Y�I@��k"$іN"�{���:��i�0�{.B��V�����\��Q��zCxT�#�':.S.]���tpuk�o�D�����ж�6�A�&�� �a��A�݉(�a�#�/�+g�+�݀Je�Q��]%�p��ٽ� H61�|����������R]ʳS�6>�d��;�����h�%����:rh�[�g*�	Iq�ip�JùGV�R#�gp��*�`1n~(�
t��<_�T\8�
i~3 �1~��1�[�$#��Ws�Tʸ���'%d��-b�n_0F!�I��UW�6�a�Vr8���y7F�j=�1>���.Z��_Z�U����ʓ��;�/�-z������D�[����5ָ)B��g5zَ���qu��r����b�u�4����pڟ��!WZt��Ѹ������P	��$�:���ה_{)���ւ��Q�5�z��gy�Uj	YVu<��E/��v�?�uɤ�1�/�g\�6ޡ�y�m���n�>�@����>i�	A3�R���nC��c����5G���\{���qH��!��7_��xF����������CSH8D����� ��q�pa b�i�JA�ȭg��g8O���Q��&��W�<���c�*�ouĮI΄����J�w�L(F�\ҿ��W	��e��e���#�)��e)U�\�6a��� ���:B��J��C���F��m�~ &Y�Yĳ��]��0@#m0�7�>~xv��@��1�ߴ����w�H|�z��g9��5���QVϛQ�{��7I���Y�r�k��?�61R#p�MWG�n��DJDh�w|�>0���SV�va�$�0��.c?�T�4S�Ēy3�����.;4}�vR<X���n�O�Q�Wܬ��P��^D�FҚNw��\�|�ߴߴ�� ��=H�ܤ:^;
�k���V�rhBͦh&���Y��I�s!yg�z��?`����*�W������٫�#KD�t��ң3k1������To��	72��8��T��dv���;}L�x�8^C��e�����{yܿǬ\�W�x��sf��j,���WP�-w�� %]���=��B"پ&��=���%b�ΪN�ԕ��ŋ/�rCt��xW��R���=g��4|e�ڈ���/Y3gTm�ѓ�1��UB�vS>�a��6��t��1�	b��F��N����0䂿�k��(�v5dҪss��K�w2Π���
�_p����6��o'���0�8�����q�IJlf\�/n����������Il2��[%A5��	�['s�ec(�	��E�*Rl=:���	�I0m����ZQ������a��J��_=�0��s�$B�#��!u~V���сK��Y]B���5	�3�^���s�`]I�y6N�Vw�������q7�g�&+�p��ve��W��}N��r'o��@I���k������:8�S�(]��l��3j�B�<��F�ϭ�\85R������2���Ǥ�6���ֳ�V�ݎj��?�`1=�1�?uf�~���W�t$mk($�;F�[+��Ĉ��/�-��ǳ~�����(!Ý��hg˪hS��C���q<_�k�q��ja2A�'�b�28`��T�i!=V�C��D��1$pcm���|+B.6�{�']��Ȫ#W�j���8�'2-_2�BW��oËj���6&�����B�1?�N�r��'�-�M��=�\�
����3�0ZgzTpB��.`ffz����
:#(��K��kx���SD�.(�V`yR�z�PWw����3��_Ç�u�ͼ�t�n�G��-ĭp����]�~%ڸ�O<%5��ߞ߆(6�*:��$O��Þ.@�~F#Ovu���Z��qyɓ�3�BC���׀��,0����V��7�-PY����L��Т*K#��ؓ��͈vL/��-�-&���\���!
��"zPZ��8L�&��Y�B�SI����L~WUۣM#��B*�'d���#���j��M�674�]ǲ��1E�+G��\�0���4������*��^	E�Q���3e\�
A��r����]@�p�� �
 :�`��d>w���w�ʟ	w`�w�R��ع���R�I�ۂc��<����<NNGI#���`[ͽ�3�-�6�M~z8������K�P��`�^��ei�9u���YO9f�d�;>w8sSo�ĕ�.��rKbעh`��+��5����j~3�oTx�R���p�890�F=��)���)낤�L/b�4U��aZ#:w��e^4y�ޚ�[��2����:� �����0:�R/�QfV�QM���R��,��UqF$���������-�8#�u�N鎻�I=��v�Yd�\��'�}{$i"���Mw��ܖjա�lh�/]�_�Iq/} M�p@z]�ԐyK5݉�B䢀��5YǾ�O����ı�j����@sS�/^E�q������_I�V�#gzw
��SǕG�]�'$�X����w�*~��b�x,Q\�����o徖g�y���0�½�/iA֒:噿_�AF�U�qH/�'�q5(���ɞj�و����׊�2��{��w�������ZO��N[���|�@��ɡ��*=��9u����ne_Xd�GV�������;9.���K=*�,j(���xp�^�D��P�,�BQ~���D��������aF�ٱ�l�X.�����B9�B�����_�3y��W۔*�fH�K8]�Ri� ̚ޅ��oӯ�U�i��GCf������� r�{[;7C��e4Lc}�'��(u�((S��6��Xl��I�I4��[�H�@E>nㄻh�Ǡ��DV����T�bo��	�V!�d9�m[�eK���DY����ۊ#-D�Ƭ�uq��v�8�TU1���D�8�aP��]�����,����%���u�Y����S����4	2�z�~���X����y��7�ʓ4�� ��������__�Kٿ�������u\���haU�/�Kg]�%�Ε��st��[P�K��䌥W��<L���(!�
/�	���$�=+w7%{0(˸��J`�wz$��[�x��m)q=}#9:p�|jd`~�]���%p+ �>���Z�b���bq[�n�aW�*�i��Ԑn�����}j�q�r�y��r�__`%�|�B}b/���C=٢^�dri���>}v��߶�͒BBc{em���8���yk4���F����d�c����(@ځ�~�RucU�\��h?3��J�W`�._��5�[?�˸t��VP3�~n�����M�
�ƿ`/D�[�'��Q��mP	��a�U�D�w6�R�gy=��r�)@Nx����� &�w+��m@Y�p���L�em����z�j� v����_B���C�������˛���V���P"8Tg�M��#�*_FH��rC��?`�荜�b�����['��u�}��q���9�Ƴe��o��:H��0i���wLN���b�MYL�M�%[���j�߬GW�n�Gß07��mf1�|x�95�����$g�jX�P���+�*��cZ�l+�b��Kc�~���̢�z��ݙj:�[E	�CM�"�J v�����6�f����f0�����b�R)س��VN`(e�� _]�|��d ��JLcY��-$z�!H2R��~�� �R��Ϣ7�~Q��YM�dr��$ZtU0X�l�"I���Ϫ8�+K=���Dī�H�d𼃨j��|ԸG�����L�"����W�-|��y*k�֡ �$��fM!:ݕ5	���ʨ�x�r�"�Ъ�^��t��,]��W���o��dk��]uY�r�O��EJ�XG�E3a:�A�9�v���J����f*؝O�.��'�������=U� X�������YB��v}LT�g�4f��c�49 V֓S~_�a+�Z���i���a3x�	Hj�;��ݕ|~�pK��'6f=~�Jb �A!vE=��s�'�U�z�e9�B����v'2��pW��lE'Ӹ+�� LY��p�o)��!4��ϐm�yS�$�������8�p�s�)c��I]Hp��ԆF?����hi?�w: �o�T.��lH^�;Va?�j<~������FsU�x�l��մ���h,VX�&�;��L�%�2lZTSpf%����2��#�+�g�w<3?7���Y�|�����1=Z���HR\s	O��	g����9�6lgj���(�ĵ�M\Փt�9h��Ya)�ğ�N�[-�-�Z�}�.S	�u�C�Y�r����qB�b�P^閰@C��F+U�7A�i��(���F������~�.�f6�tI	[�Z��;�r�� �d���^� a6�$�����o����"k��P�2̊0���{⥌ ���8�Cص),�����f/���^Rq������eE@���yRϡ�t�1�]��(��{5l����oR��}^��428��;Fq�@y��A���}�J�$>m�]?�un����x���>���v��^D��ҩ?{�K�e�1R��{�g����y􋊠5�\�dGfd]���C ~��š��f(��*�,0�fޡh{p��*R���d�&ə�����A����Jw�+�[~�
0�qn�<k~��I�uGUpH����'ְ_��o!��C(�J;Вӣ´B��}���a�4U��0�!#/=��C#-.\/*�.�E(L�鑘�/1KN�ú"�a�;#��|�_�l*q�|��ܮ�0�_���d��j��`P�e2c�O�9j���E�XӐ p��c˿eQ�DA��,��L�~+*Z�G���͇�Zv;�´AdՏ�[�8�}Ծ���4��6�����v�Q
@�R��cza�˺Q�.}��f2�a^�[�$I��DC�/����hB�]'����U ��<f"��%'�w�{+���.u�kI��0��Ņ�=fh���<�Q_\�Jt�����'�:�Kcʈ�hǠ��9|��o�r��Į��z�t�ۡ��.�	�}�NA��Y2��[o}�j��b�"�xXYH��xX@ً\K19��ވ��D�<	��J�,�"��
7i�� �ix�c�
��Pr��=�����V���9��0��J ྖ��!�J)RW'H� �sc���~�9�V��gᤀ�"O?:)pz��"P�M���/a·&��
���	<�m�\Ҝ�4#�P��}�竷-��3��[�t��?�]ҘY��)v0 �K�������V��uP�</�'�������?�]<�B�jG�C�����k����a'�e2�Ã�۶J$wf	&�3hI<��&z��\�G�F��[�fw9W��r�q�w*���TA-����V�(mM�r�<Q�ô�a9�E��Gc�;TcpQA7W��:HS�r��W���������%�����T�F"m��5Z�i�ڹ�4��!��Һ'������Ҁ�5�FW����p��۾�:�q��^٥&�u�\�+
[�o����&*�o��m|��X�Y�n���\J�)�I��/Lk��qqs��I ���È�^�L�yfR��ȕ���,�&�6v��� <`�ɩ=�?t��DP8 P��=�s(��x�A�I
������N�"7���xԕ�25�w8�����(k�P��'�?Z�3`6-��Z�ѓ�^u.T�2m��h���ZX�3���g���΄\�<�0���R�4$8pڵ̓�zoC[�7.W�'i<�P�7� �;�_�=�7pQ��>�x��[i�ҪN:?�
�j�d$��[&�,#�-��#R#��$����a���[Ʀ�Q�Q":w7�i��58!�q�}����4|���戢χ�*����JG|�W?&����w�.N�w�z�MQG�=q�L���Kh��'��5�����	(��`�|O����b ������h֪5�kj��ڙC�#�H*����l�p?)v���{az�vҊ�"�G�q:Ϥj�U�)��⮺����g\ٿ?0<#�^�au3�np�7ANM�?�`��"�w8�Ox�b� pt׻yi8�j>`�pYHr֠!1_�����ekɇ�����]CV�c�i�t�����K]�7�@�9h�gξ�6lW�&�M����O�`E�����8mR���/Z�lMW��gcO�y�W��v���D�|���g�*(����b?X�U����o���K�jjG�m�m�r������a�Xz^��=&Ǉ��r�v�uXBG�	w��B���4��^]l�V�l�}D�:�򫖩���@�M�^�n���`~�n��˯�6���g�Gkv���J��c3�g���2*%�3ޒd)0Ϟ{.!Sre��@��q��/
�
����-�tè��T`µ
��G��`����L�):Z��*6�����I
�hUQ���BG�H�XA�C���n��];XV7���)�L+���XI�1/xR�2�h򖅫/���[�Fʣ��;�i=��Et�D��{����Z��p�
3B�)��(����=mK��~���{��<^�f��Y+%С����}�b �I|�_	"rc(�R������)e��1�K�>LX*�W��� �,�{�a�����a��߀4 �+s�3�ˀA��{wҲ�Ow���L��R��Lt*Gy�![�� �7����&���~#X��[��Tm��XCx��i-��c�O�Yv�b���Ն�	�'��?�K��+�VF�t��;�.2�N[��I,�_v��`�-�	��ag􆱐�!,��J'����Y�c���4&�O�mU�l����DDP����&���ND6oUR>S݉,�ό�jYX�Zg!9��'�O��@38kY,�gGk�c�<��ܠ��đ��/Ce�=��5B7%�Gs}u�'f�F8,�t,�M1H�B����)�@�jũ�Ώ�>,1�$�M�l=���g��N˜޵�*�>����(����C��թ�_�&����&V����4+H<�.�^˓+v��(\aK4�v��GM��_�A�D��d*LCf���ҵ�\dǯ��ZUs��Ur/����c}��&[܃���1�����AY���O������kw�]���	l�����G���}[b�GkGȍ��g4fk<�S�M�I�ﬗ�SwJ��Vz�����z
R�����bG�L Bڡ�gH��������ҺKWj��wHH<���>�X����`Ek�|4>��XM��@Pj��8��ԅ�+���{쀲SdcU�������j����ڔm���)g̿�.1W���1L	f)-\ωlZP=2�1�nA�K���<ͻ�rQ�
KuZ\/i�!ww����+O�=/���4�5��%%�4�"�g���F1��0�Hw|A���=�Fӧ��YT�{c@�ϥ�y�+�r��""$���T�0�p��|�e�H��}���P8'U���l�"���րa��g>�^�Q�.j)?7�������@f�G8]a���W��y�/��{��9����ªs�00��r�uqk���ڇ�z.���o�����#���x�Tb������e��$6wЁ���m���m[���;w��X��������4��1�(�fVڐvCN���=� ��[��~��~!N�Ze	z����j��ܑ_����������cM����Ӄ�u���x����ǰSs�.���C߹%(.3۫��Lpҵ��0�2!�5ol"��t>"��F�����r+>0R��	�7&��+����W��s�� Q�<��K4�W Y���>��2�^�g�RZ��@i)�f�dH���`?�� a���)VWF~��U�7�]�<'5��|+�2�D��T�G͝�42�ugT�fx�����L���O�� ֔�3�D?'��By.�&u�.ZɝqOٗ�/h��ZX���֤�����ԙį�X��%-w��
�p�?g�=B������~a_�V'�Ef���*�WU��@�N�S$�~�s�j��4D?��B{J��R��[�?(����UⲐ��%�r3
����ɻ� �tƉ@�`��*s{tW(9X.{�u+�֘{z"�O-�f���qԎ��w��~S��ܱztY���W�K0��#�6�@�8sb�w�/�e�;u��M��K¦���F>���Q�t�}� W�S��W�\j��,�4��C�a���]e}�1�Q8��IGۄ����f�N8z�P�䓯0���Pvjƍ������4�-��zd�����ݔх�ʩ�uY�1�x�x�J�Oyu�y�ZV��X3�|Ox?�\jo_�ȃ��1����Z��U}�ax�ѯmZ��
=�^�$�~Siv�0��o��%�2���d��.��ܽ�%w��U��8S�%a~L(1(#��6"i!�@�o������������'o��� Q�!����/�j����s/�(4�ֳ��fD7��sD��{,�&�6򙓊v�T�k6Gi���&���羵�,岧+|�_�d9��3�u"�Z� ��l�~^����ШT��f-qi�k��Lw\�n�7��PT�5��%�����3�{0.~�wDc�2���"ަ�Z,�'�oX�^w� >�|��}k�#Q��+�n
�t�
7���o�o��X� �����Nd�-�8A#��i%d�����*y>�p�ƇC1ڈ�1�k��0l�x�J��pC�wF�t�#���=t�n)wu������ 3rI��G��\���0b��_f�N�4�����ߗ��䝜�X�w��g+��W��q��x#�n�V�)�%���(V�&&:c
�6\l�ؑK��S!{�����H���;����zO��p�8�T^>488:�*����G�ʨ�M��,�\R�}�1�R�C$u\E�҂�bx�N8����24%�9t��]�����Qg��(=�6��s�_��G��7��^[Sr�9iiu�xd����H���A�I^�)�Vb�lZ�j��_Y��6M"�|�ic��ejʢ@�w �s���o\]��{�*v��RS))f�<sn2W��c4�73=�2s)�]���i�|񯻸�1:��*�.Ꭵ�YP����iX9a���/"~ ���z�ϖ)'���޾qU:�Cecyg�dJ��K,�ֵ[��]̖F�_����ߜ���g�#	p�i���T������PJ��\�h��壃��}�N=�e1�w�X���͑�,�[���%�*�@����t���J��T�l/��)��B�pʬ MY�U�R@ƨD�_�
>��A��Q�?�82
��<>���v%�!�S+�{�'�]'�|�T!Ԧ]>-�1x����<s#t�+�[FL}N[�5N�"���+�\�����<�4r Ws!�d�u��@6���`!���j�T0����
���o� ��n������~��H�v��Y���)���o����鳬���H�q�6z�snO[��d���`�?H�)�=���;Oz�Q��ר;�af��|����p�EN?*����P
q��ս��������s���v/����ض�vx�@E�RD�se�g,<��=�=\��tX߭��" ������
jf�5�8�� W�}��e�S�O�%�����$ٰ#�Z[.�U�~JqÄ����
{��.Xs�;�9��E�\9��2[��A��%��c!�2��-o�/�Fo�=���S̍����+Tr���]�Ќ�"앁I�:��4v9<����v�yx��υ/��5�yR�d+VtR��J��/i����?��{s�=D��vGap��cɴ�|N_J��6�U���Ηq�]��ȱWj�"�y��,�ƚc�]Ð�:�����"�eu1���hB:U^����Pt0X-��\��ұ!�F��-��f�]�5Dc��_8��_�����˽�C�̖,k3�Yz={�eP>��U�y�7����]�_�kJX��1b��P�k:"��`��a���h;�b�+,��f-K�T)��9tt�镕T�aG�^���H/g����J6��M��a��,��u��{�BE��2]�k�)D��=,���П$�#h�)q,_���C�Pp+Ӿ}!p��4KΟMƪ}\'��w�v�qyW� {B��2�@s��Z������pa���)��'�/P�d������M�~)�	���l�%�<�qy�[�M<�xEđ.���֌��^V��U�gi]�Ϫ3��u���S�*�8�L��٫]�aTԆ��-�� �6��Rk�{�U̜U��;�V��szd���wP�����m'N���}J�<���a	}7��0����9����ӕ2�?A�;��na��=`pW$�R�}��]#/��H�3~{��w]n8�pk�)��Q��h�ZS��N������+\�����������*��m8
DZ�]�\9Ɍ ����S�٪
辔����܁���)~�H��N���������������/����mm#y�����I�#�^Q�:�"f�C���t��e$$$�:Ox�|�c*B(���Mc��V ��)ہ��7~	��0��A�wFyL߽růH	��h`]�;�_�F�i��H����=���ߒTjK����w�:/�a93{/s�!��2	����kS��jhJ�[�,ݸrx������gs5����f)=w� [6m3x�|Y!����w�W�ĚS
�kr��4�����������Z���b:�c��Qv�^5(��r�}�  |���r�i)��P�,kF���S�Q��eC�m�68&��da}Tѡ�F5�t'�m��b�s�G��^T��K���,NHI�|����wZ�;IN$؋�CD(:3E8`�����+d����h�a!	�r�ɎD2O�~������I�ْ���F�M���o�ʇb�>�U���d�������N���Z���vZ;�	Ҽt�.�,��3a�������*�:�g����R~���Q� 0uT _Y���	C>aTb�O�A1"QH��i]V�׿n.L� ��3�h��B�oC��i����$����<?��U�瞖�����&i�崽�:�yF�S�{˽Wc�� �9��8���j� %αi�yvfn�e��J�I���2�Av�����.W��Lv誘E��v��S�sOd��
�JD|�.�y���9��;"Q�ߒ6��񸐣.-<3�%�SY�a��r���v���U��(���e�0����M�G�E�Ou�V�O�y��
�Dx��)����%V]xAn3�@�~V`Ϙ�#z�I�����i�#'M��gw|���j���K�*�_8I�sbd�6�,�x��y����ee&���p�)���'��"���` m5HŎ��Pv��\�x�?n�k�fq�_�=��'9QH�/�\L�O�؛�_�n{�̙���3�	�b�_Q�"trO�$\��
�5V��9Z�l�+>!6�ț�k����c�p�p ���/�e�wn(]�����S$���q>d4�j�HN��)���RC}�B����z4�L�0�ǖ�������r�7�1����'��O���M��K�q�k<U�'��4�^�� �Yza�.�4T?	�](�h�1#v���U�p&͠�h�xn_����Oç���,�tw����c[�S��!=�2W/�^�{DX��_�j���[���\OR��몠��K��WwD�e� i�N��3*��u2�-p�a�}WtZ��ϜCxݕ���gOZ��@T���3��.B3�1�D�[�i���)�� &t�_h����mv����/��f�?�t�6@Y����e���1��s:\�ǂ�v�e���o�\?�U#W��T�C�Z � �	JG�YH���� ���ǯ����{8`� s��R����[c#~�� ��PrHsyÏ��l�gH	��)'=	O�7�k�C�m���8�Q&�/݋i@�g���[|����xyh��|s˽�ǘ�L�����`��Ư�ai���7��HZ	R �ܰv�s�
3�$'J�%8�*���G�GB��id�?�Y��<���t�߇��x��9_��moz�&!	3���3���� ?@���e'�E�U��+��x׍!'?�)?���iޢh��"9����
'�cI���<I+��Y��V=$J���i�&�lײ+�/�)͉6Yل� ����C��qi>��|"�h$���<���B!��/�T.-#1�6��IN0��j��eְ=H,��K\t�!��p���Jz�Р�[�#����0�e���HS��ǔ�ĕ��a�T��NT[�K�n��~cU�W�8)�+A����Tv���D#Y��V6ĺ��N��"Z̻��~�\Ÿv`p�3����ct��0?�r�ǣ'�"�#�,��}���%=���"� �K͙;-���4&w�sO��J�n��K��ژP�Lq�T�jq�a-n���<J����|�*/�N�i�����R�Q �/�c���w���7��N:�7�ޅ����.^&��Ɩs!]`/�f�G�4�<3;9���:%_�GS�5j�yo��~Y�d����J�y�ƉBqf"����	�I���2�����������u���=�ړCZ�Y�qʦ3����=ٻ4�w�;���.������-Zp�<�BHQ�z埬�V6�����{Lw���]������orO#�ұڷ�<�o^��Ή���F�7*�hN�L����K�]�J�|��NU��_*��)�p��ci�Kd+�E#�&�N����A����?�&s��a�s�{�0��aI�Μp^+3�3��o����WH�>i#�ރ]����m٦L�>"���g�
32�Dv�١�����S2k�5��|hFٳ$����gL������Z��T�l0�v��A���("���2u���BPؼ[��!�C�W5�S;�}!�'��̡9�XvQ�g��_�-T��+`��"�e�w�$2  3?��3/CF!v�S���@��}�d� L�y���x� ��0��Q�&�8|��������kRR�g�|5�<� A�����s���b�������1C�3�����Dm���ڙ����"�R(��Zu�A����e9������6�W��ً�c�xZI���@&�TQ "9�/Ur'�؂��GxO���<����N�<�)��t�?�~.pL(*�aS��`�£�5-9�r�^��:xy���F�5�L\}&��z��|V������n)o��n�3ܣ7����c���,u�(fF(2��`�7$�/Vm�W�v�+,9��G�;r4�-a��*�*�s�� M��X,�6�g/��f|{oou�̶�v�W�Ã��	鳝�O��_k�8�EO��U<��J�OM��:.n�Ő��G�f����"��
Ȇd~�/�f�#CJ�L�e�w$�įPZ�ڟ�q
d�]b��6�ݯW��.�>]�C���n4�Z�V���4�1��	��ܳ	T���?�Q�*�X��-a\�nI`�Wp�1�׊ZS9�8W%�R�ջ7�w�e�)E�VMt�N7`[0lAV��U���!��_Q`��U���cK�@
�B?͓T�Z!v8�@�i�ql2'�͹��$m�h�.hΨڷ��*�E��_�Z	�xy{��z��u��ߌH�]>,�i����L
fC���g��8�$Z�<Y1Z�B!x�U����b�f�S�0J��m*���`�-�O}��y��<��g���>��R��ȇ����˽��IV�x��䒼a^�[�'[�1ú�Ϻ�G���3?!h���?OZ��_]�BB���� ~�n����Zw���o���\h���|�22̴�{Uw4�Ⱥ]6��+��װO3�����i@nOS
EX��lř�)���}�ꭢZ���F:����kL<�B�0M/����h��Pq���/EV}����nZ���zj�ND�@Ʒ2k�����G�Mdε��1|�~�H��n4�0՝�3��gب�5�0��Z�w�\�H.6(��V�툄sX�Z���v)s;��g<2��� p<�x��S��:��~}l,�����jQ����O0,�4K+X7ش�w�@pJ�??Hi��w�1�%��Ζ%���׼�#Tf��A�H��=��/�g�S�t#�`�F�И0v�cx?׾���t��[�M%Y4��e�P�t�)r���TSK6Pr����0�?V��L����s�ұ�x)dw�kF=��g�����WVjyn_y����+lJ��C��a+�[=�#~�\|��E�A ��C)���[�'�	�*�G�mSz��:B]���	Q��a6�C@���p�\��lO��>� Cۢb�<2��Z:��4f�ʙ�2S��6�|D�{��l�P�������Y�������L��u6N���>"�G��H��+��K�#ׯ6k^) �Z]k\�w6f��)���.��L_���T����jL\a`!��A����7*����Tz_[KT?	�:��̖�I���%�X��c*&��C@��A^�z��'bk�*�K�؞�w.ƥ?��x�t4����` �I7�+�KK7�rw&(g���$J� �>�F��d,.DIq}�9�'�Xd%t$��4�q�����.CbjJE\\薙Վ��tR���I�+l�a��##�E��>��gm����4�RL)p���ڭd������$GGhY�o��X9��N�E|�4(�D=Y�PX�6%,�h(�V�����c���%�nq�&C6�0Z�1�(��ў�G��	H��4���T3���I�7�7�!	Ĕ�}���|h|��Yba1�b������!�*�ƃ;��^8�'ȸy�T����-{Z�<r#���r�u·��~B:���^ޯ�j��a���P���{��m�o6R��r0��~�A�K�6���CDk�0T�!Ⱦ(������zڇ�v��ma�4)�^dׄĐ����P�-E!����%��	3�g��+F��r�;�4�k>Iї��&�+C��t��~���9b��ʊ�#sn�Xt?Q����9�赖bFS�-ŵa?��q���i mN<���3���\X�)��f���d��ܞ�؃qw�V��W���ܛ`��7���73ﮍ�yHs$Џ��������ۼ��(F���������� AR�l�lS�RǪ:A�R��%Y��r�3�X�NI«[TAԻ����) v���o#zK��S�=�d'_�s���B��\\�@�"���Y�^���@�T5Ѡ��2����(IC`VFk���uc�4�q���O�?�[�'��G�?��?**��J�Q q��6��4a2�h��fv�*hl����+�Yg9e��X���B���=:��Ɲ������r���D�!d�'�C��Š�_����?�>�5v8�I���d�<�e��U�)�L|� ��9��g�:��f�����a�7�Q�H!�)oE3|���f��D��"%�r}!6�Y[�2�90��8߭nY�J�(�~mL��b÷F�����.���L�;ǘ�����}�2:B�U �_�Jb��͐�h"tV�[N�78�p-���Z|�I,f�~��)@��"Tc)�aL@��+���U��1@Kk�B���u��o.�����9��6��M�,k�nd^V�t�@ӫva�Z�T���ZZ�����x�f�T��-服8�FΟ���El���nlK����I���B����4N�
C�����I`1tg��Z�{�m�0��P{V�����.�J>�1��L��{c��~���cq�Evdn�r�tl��:9QO!Q��g#�M���͎A��>�ge��L�E,�%+�y�_�l8�ۮ�7[x�m�0�;ϧ�.�g�m�h�F�	*Z2�h���`q�W�Kk3�/���,��}.-����O�K�Xj�>}�MU��lk���\g�X�7��elS�t0��Ϸ$���k���F�@��L���M��x�I�}��H��rʗ�B34P�f�]��Oc�)Œ*]��h0�� v��h����ї��Gr�
����JOW�S�a������}���Q�@�ˣl�����v� �P.Ɇ{n6ս���bé�����'���tN�yb�%��p�p�I���w)�!'��	�
gA?��jc�鳟����5�O�i������^U��)"U���@��"'&�����2mk��V����lQql�(d�K����,����~���W��+<�rm��n��� �MK����=4��HEFaՠx�f㴹$*���:��Ww��d֦|�*���R'�	�V�֙�T7��5Zǹ���+�8E�T������ܭ񝎰�!���*���N~jM,��4Z,݅7�K(�º!wf�A����e�c�db���$���gf�L40��Lo���F`�U>��D�M������tmF��bTY��<������0+����T��c?W�T��{��pn��@��z�b���;� �7Х����rIJ��� `Bb�,�<�����r���P�t��KZ��c��l��p��xܓ��*�w����γ`�"d��#b����o�b��-��9��W�}�0�<v��-��#�(j\e������o]>̐�4h9�@�â�*�֘���e�Sg{��B�8>��*���r��AN,���%4��8n#��ύ����5��WR%�����;D�K��gJ�)�<FR��5�+eނj���`|kN(�o�z����V�L��-���{z.��}� U��������L9���G���(X����)�v��(� ���xmTC����G��tgD\�<�j;���~��ֹ��Q_f�Q����p�]-ߥ1
nQ����@��;�����Kȟ?-�OІE )�����k�Z�!
`��֑E��d{�*�1���TW<b}Tx��I��r��H\��x�Y�*{����X��"+�OE����ޑ=��?Hlʺt]�0ux�� U1	jv|�;�K�O�ĥ�@#U��H��+��I#��P;�دL�H���Ճ�(:��Ĭ�:����=j��&b�U��F���3�_ֽi�{w	BY؉�T>2�萣�B���B��E��u~��(� L��Fy��%�&_����*]�b)���l�a�X���UUF��`m�6�G��V�}�B!�Sj l	\������GP�  �ÃgɌ���/B3:V���T�u�ל#*w��a�i�W�<	G��x��T�Ӗ?�w9H�QC����({:��ק[l����G����v��6�;�z�4TN��tכ��$�_E����<��+��X
U_=Q�0��3�y-�RF�����^�"���S�N�vq=G�2-2 &��Hn:���f�Ť���Q.�d�������	{a�uhv�i�0�z(��B�&����?�!x�q��h0x��V�Թp� 	0��m177gB	���Gb�nk���턢�m�X_g��=��!QV�
;��x*6�葺�h� ;��iog��l������]"����-�>k�}��UPzu��c��eyY䃔s��bZ;u���V�'TL� U%������-D����$IZJ&���D 7��(���8���]�����"y�l:�]P[=�eQ*"g(}ʔ�Y6�"��O��&�6(OPD��xRQA�$n�,w`|�	Ź3(���⽍���%q�3�� ���$�`/���%���oK̠c!�+\ ���	���s�_X�;�'�Z�ݐKL�N���ԧ&��Z�e�ء0S9)",I��bǊZ���Р
%Lk��LA��ͱ>%���N�reD������\�x�`��q����
[��xE�ˎ�9��d��~�5�D��"�.��8�9�iC/.�v�b2�g`D��v
B�$HsӍ�Z�/��)��j,|89d"��O��OW��Z����֚��H��N�$4����:�1�3(Ħ;���x{���(�u�c|�vT�&�@ ������L��BK�=O�u����M+���B�S����f��]5��Y�q��cIeO=��s��\ �=P1l+s�V����S�4�&jV�JĘ�0��F�p��/nÊ���}���O��1�0j�VFB��9�w~�n�<y���ݘ��j[p2�PuSK�����rH�ΤME�|γC��ǡz�eơW�v�3�u� }A����@�$����o� �Mi�;6�&�N+�+G�d���'��@@p�u��R20�i/g�1t�E���c��r+A��F��T}�;�p;I;)�?t����W��_�:�Ea���߼��w�u�m��w�x�%H�	vIz)�n�A<�!��b!��6i�ĳYS�K|�\��P�C%0���	�7y2�z�vH`:��~1P����b_�I!�A�8�L��A'�J�O�	�*^�S-hI�<�� ��xP�<R�8�*�8�¡���T��v9MW����<oQ:��^L`�~ޡo`</���?]8�~���)?W%ҚVP*P��:�zu�h�!~��qכ'�������Q��[��,�P�
���խV(��)��VS�oz��?F,�.�lw~:].6Z>�]��r>�I�V��h����ηq����yY!G����r ,k�%F$�K�|9��/���.s�^q���y�]��Eެ^��m̞Ne!zG�.?��?�)D@��(�Z�wf4|:YP&3�!L�5j�+�y2(��>#0���Ѐ�U���wE���{$��ȈM鹛�E����xe[z�������Ď�4�j��Lܸ.�ۯ��V�A3�&�$��_�Ź�Q��V|3�CN��K��~XwB��W!�j��	k*n6��X�"+~ן��$Ȏ��zgx�l(2�I^�ȣ2�5�ÜK�U�tA��mr�5���7��6�0G	���K��ʄ���L)}kC�qSg���dա��������\hwQ�w
�h$�����?��?�<�24��Rc(��&���|a"�*\i��fK�/���<��9�:#�Ȇ�5D���C��g�ڲ�ww��Y�����k�q-N!���/3��ޓ����G�O��P�"��sT ��/����Ni�H��4>n�9��@y�S�.�~�g@��6�n�JܻMsl�R�i�s4S��̜�}J�<<�!��yuu�Dg�b,�7�Ԩ��������l��M0M`���/��h�|�!�������S�|�s����ԺuD/a�)T�Cʍ��݀�?v|����HM���00E٤�b;��Y�X�ty��d��7^�<8��2�Ԕ��:�v#d���;A�B�Tf���2:���x��QZ���$�g�%'#�~�˳0�;�~�$c���4k�5r��y��m*$FkzM�/FQ�	�5F� 1��k��\K�Ț�(�N�N�--�ŵ�!�k�ywR�l��ޑ�$+�	�n38V�j]���������)� ���=C4ջ�?�^�<L~4��v�lx|1�"�%�e���[�;���P�dpߌN�������~
�0�x�܈w��8EQ��+v���ȅ�i�z�x0�!p��z.Bs��H+��y�����`�^�K����l�������/%��DL��K.agN�+�zE���S'�P�9���s�n�[��)3�>�-���H��m���������-�ۀ�ΫnW���K��d/����,���d{a����05'0Z��
sw&�D�t��-z����I@��a+�����<?�vL�gLO1��)^z����Ҥ��t��wB�}bc/��{�h����;�P��Z�5���u����c�4�H�l"5���J �|1��e9W�SOڊ1�2���ED�σ=9`��Q�f�WS�[ʟE�k��j_��Z�qБ�L�Ƴ�) 6����X���9�a�Zwj���J�X���rO�r�լ�E{g�sN�ࠪ
t�?@	'�8m��h��eB[�]�\B���@�}��/��R��n'�P��!Er��b�,u��D���F�q�0�*�|�9����C�y�x���u:��${\���SƷ����p���я�ú@~�d�ts����1r���9�;�興�����C�츂B������"M�}>x��q�,�:�V<nf�N�8=a�3�$PV���Y��2̧���/�5uX��oVz�7u5B���}���	Q*�{6G\��/oR��y �ЦۂI��sqg��!�G�c�q�sa�������YI�����K���:�������Fn�_|ʃ��;���PS��L1��@$��n����6S���x��f!2�_x����G��4~�kq�+�(���#�܁������_��MB�i��OI�ZP4+�DM�Y��^�ypeR��!!%{
�%����8�i.	5S�1�K����O*���pX<�$n
R�H|���Q��_S�n�qmUM�G����M�iI�%�iK2�+`�Biy��/�꿘\��t�<Vl��?���]��;�4�%=��)ܼ<�ȑ�r�ұP	A�~�,�XrA=@����g7���!��3\���֣�'7&d���)�@b����	%'*�� $x���D��S����m"�!�ʟ�|!Pf�^w{㻊�i�(���3I��=KђgC)��U��!Uq*�"8dA=�gD��w��w��,�P%(+'��\�}����3,�6S�Bɧ􌱽U��5����4VJ�����Z��5���,4�v��sc�QPC�,|f���Q����7���9���>[��爚��z�m$����/f�{��ۭ��Kу�K�qQB.�8����U9l�!���W�~����jA��>B���+]0+��Ua�*Bg��������1��Q�Zvv�l*9uSc�t:��;�`")#ֲX�~�/<,�<Ӟ���F���ٸS	���E r�vc�d�}��q���{����"=H�{܁~�]�=@	V�!�J��}�������э̀�h*�Q���v�x�-�@L�^\#떙��T��Lӱ��������j�f~��*I.KȽQ2T�1h�	���]�!$e~�>a�6"��/R>\8\�ok ���n�^0q�\P7�S���@������[�d�1��$� X�v$�R�����zHHILJ͒�`�����r�M�[&���Ґ�Q��~��y��H���Ҧ��q�OC�u�DYt�3 �C� ��33��v�A[�}��僈;,#�U��ƌh�5���8�3�B^�j�V����M�Aϒ?>���G����@�]S���U�Hև",��,_^9��=�����!�9K��
XKW'↚�'oid~��T������\���6>��ff��W�k�>7�W��0�/+Sz,���t��^XGؘ�xÔXk�pJ�T�7|�Ϛȍ�u�ؐ��ԔQ����y�<�����n��m���t}�:�ƶL�U�Wx�eLC�gO)�.:;-�S�� �%f��L�[�ѾQ�~b������>�r��s�g�ŕ�eۊ�Lֱ�~�eĉ�����3t��E?E��B>��R��f=.��_����H_��[����i͢fJ��%��1�5�4���f�?o�x/��c~{:Y0=�?�ԥ	q������v�m�}�a�.�������_l����q���a�� ��61�E����,mꕁ��h���u��6�S���u;�x(7�L�yL���Ͽ�!��]`�Y���L�|)SK0Do��?���3�}�m��u,�ʧ����f������y��E��O͜Nɋe�;�($���C:�*����z�b���ٶO��)��{��|�6�yk��ћU�m���̀��$F�\c�0���,����c¨�K�Ȏ��m� eY�X��4��r$T
�%b���v�;k�o|��&R�g��.VGȘh~U㓪���~1(5M�"��R�OҞ��{c�V�����hX*�Y3�3�BP��>J_w:s�/ݪ��SF1OYS�P:W)��)v�0�R�g�Tm@�w'����&�m`�R�4 	��2ӣ�.�fZ����l� W�K���$\d͍l�M^�� b�%��Y�/������4��iF��om4��&��U������M�x�^��$�]����b��: �R���	.���m��<?�-?.�rtd�!���U�H/��?,�,�_��U�����^��Ho���)�C�GSV19��j\J���l�ȧ�ָ�+�f���΢��;	����͘��r?Jʌ�ɮ�c�")X���)��:c!��¢V@��X`Jc	7I�0� gQ�.Ő=б��l!� �����#�_.frX��́%��E�8�^�d���U��6��վ��^'���Q�	�a��g�5�#�;��~�r�x�LT�=4�>�t����_�i|����^�ɻ,L*Thv.A�Em@�i�)yY"�8L�<�j���6Zv��E�\����9NW��É�� ��hU���Ϳi,r$��_�ì�����^�ց��X�n�+GJ��k�`��Te�h�B>Z�1���R��N6��Y��Y�$0��?��!<g8��s&�MH*���<��D�&^>�L;ң5�[�y���1 #��6�OmO��?���.�]��mC;�#w�����#�#�F�*Q�L� �V;6j�u����!�V���z�`~�iYb	.���;J����vJ�׺����6=�^�&rZ���}�}�b#_����?��0sp��0�T ����(�Q�h�$Qw��q��obʑ���2��Z;̒��
����=�X=F�M�щ��jW9�EU��D�N-����C���ɩ�l�%��t\��b{�����/�9/�i	�y���ݐ�o����	ɫ�P(�x�J_� ���`1#�^�.�����7Y�(
0��!�/�f����z,B\ �_�k�2���l(��o�m����;Tp���
	e��n�'U���aN�(<��=^2�ȑEl�y6����Ġ����db���*X&�X$����!Z���{���6U�O��f��N��އ�B�ĸn*)���kmyUH�����_L��]�=!�����y���Cy�m��kE��Iؤ�[m~2�*�W�:v��W���Tp@>�#�c��nA��@	�q&�2��0#_�% h�C�I��/T�8\�<�3m,���0-(a��TB7����%�i���kh�1+QV���N��;a� ֠���@P࣠ck x�DB�<%�9�tN�p��:�۞g/�Ť^�������7⤱�U[�V��^�ܻz��4���K�&ڒ)����Gx�Wf�r$h�5sq9��?�ĿS$�GM�/���>��������mJ2�� Xnf�F�I�9�!������P>�S ��u?�Ms�z��1�vm��s�L�g %�DN��9�M���D��ֶ�N���+���V��C4�2�Y*�~�N
��d�z�	��t���#��{.�.�n�^ϮB�$����q�����~��<������8��G�eܒ�i��Ə� >�p�� �o[���[��CGQN��]u�s1��/3�*��x�Jʄ�(*��╆�)���^̢V{E{i����9gro O��\&q��9f���3fDa3� �˷��{S��<�Q�����U9T���7Zh��M_�.��i����b��c
 x�Nu?��fϣ�,䎦	��u�O��d���k !��h�b��E.@� �A��U/p9ܛ�7��3�]���Vz�V��B�G���Y Q��TM�fp����$�j_^X���7�&�Af�Q5��ϩ�#���ֶ�����w��pD�\Q�f���Pl�}�*n���t!ֳ􅖘w	B�ia��/��{���!,����,I�޻�	����p�R�ГJ�Z	 0w|^@h;&���7�%����P"�2��5��"wq�s�t�g�p�"A;�j���+C媥�Z�/�ί������t�D��f/3:�%\ː48�@��lH2�D"n�t��2Uz}��p�YA�D��y7o=�i��ma�RBQ�c>��b�"+\�o�n�"$v��Ӎ�[j�G/�;}�y"��*0]����<��թ�)���\��9�NNJ����)�E!�u] \��9;�e=*���`�u�#v(#�+:�8��F��ԇ�1�����C����6��7��U���3N��N��>�W}�$n�H���}ń��i�Y���Z*ʙ�#�� ���e_��=B)�>W�C�԰���6�`�"rH�bM�>a���7�F�eR=6e�dG�E��7wr9��q�$�m���	�	���Õ�]�j鶰U�S�y��k�LaW��s���:�q�.p,���$�K�/���7Ε�?�f��A.�k�e�ڻw�?��C�&�7ȺR�eQ4�9�*�d��Y�C|Ӿ&UGl���&l�g�pU�V������L�_c��5��t�"0|�͐�R��,�Q`��g�_.2����乚+�o#JERϔɈ)t�F!ZU}�yz�ߐ��pLJK��].WX��E'��9q�}h���Gw3|��h Z���rhT�<�?�o��Q]�qO%rkl/��-=g`�-�?6�ۓ4F�Xrb���όlI��Ԫ(
�=�+?�T��]P�JT`8�obN�m��!�"��i����	�D�!�vl��x���|�,:�%.���A0!��k�[Es �-0 �5!�	�v��	ԩR���
�Y��������ɪ4��d
d4D"�vf],�A��cv��&G��{�m\�H|*tb�P`Z�e$K���s���_�Wf3�[���Ŋ��U��+L�?�Yf�i���	#!�!$ܨHa�JQ�%~����T��+!r�]�!���<+,���V�K%��P�@�>��v�t���!AV�Ov�is���y���\@tD���l�{wE I�O{'&k�:�d�w��hQwڋf(P�!��I��O���M��p+�Ӷ�c�6������-6|����ڔ0���;d�X�AA��Hv���2�*R�-BeKC�7B��1/]�<�B�l�2b�f3u���� �&ă-t�3�?���u��R���p�4���Q��,��_��ah���ߝ	?��t��z���L�S��$�I����a�b��]8ta��d����e�Zr�nޔ�NiE����6f�U�=�[ ��v�X�3������hU�[95x���������M�K�.�y؅v4Z��`��Y0J�~\A�KI�\���G!#ѹ&o�ң�)��>r�Q?q�\ʁ����Sd�,�	��U�\+���gr<���0>b��/�#��{�]%�I{;�r>F��z���s�\��P��Ҳ�9�79)��yrz߬;�'l��*��X�Tb+0�#W0��U`����VR�A2_�>�J���vu�UQ�x{�U8�\��nHh��\,�VD9@:zS����G� !��j�����t�7i��R��}��g�d1��+/�5L�U���`�qT�>�5�#j��aiz3A�磛�ﲂ�b��(@z��E3TZ������"J<�XJf:��P�!$�7#c����ƱRzO��7���a~�\K���Uk���1��YV�k���v�Q��ߔ�2��<A葪�Q�\���"mTW�=�aZ,H^UWB��8��]E�����׺��lo��(&APe�������RH׽nlEV�+Җ�U�(���	�x�,�k>��[[Ц��J���OjF�F}�ѭ=;r3��SM���� |i��L�@�����J���W�3�6�%�6,NUEg?<W"J����m�P���(����؎�e��Z��M�� �۫�b���y1��<+N(��!8Y֋�D­]���e����1+�g�.�}g��e�$��[Ȍ�
ܸt�#'Z�+�9ƍ��#�S/4[`;�u8u�,���)��������^P̀"������#����bՓ���g�%j	�Xg��/h�|o���R����՗��(���] 7M�7}I4]C�K����O�Ε�(֋�P��H�Csa�/�h�LV:�W�m�8�0/xԀ�W�NOpT Jz��\���Mk�4���oJ3����X��c�����+�����V�֟��ڌ�~�J&0D'J��Lƭ��2p%KVM���*#�L�n�Ľ���'����e]c����G�pE�h>��>��	3�`ހ������x��m�iq��U�o�>SeY���8��I�<O��7�}�v���7��~��S���!�B�������U͡K��%Ý����ٽ�"��PZ��m���}��Nd�Sc�,!���Ͱ��,OB�u���g����yeУ���2�w_�$�ْ~h]��'ym51F"����ق�� "�}1V�M���=u���~����.���]��4��h'�|�K�h�&Ĕm§��\1�w#c�n�Y�7bvNԅpN �v�֦��8J/ͨ���I�		`��9 \ޠe6��P�pJ_��͙o��;�Hx(�4�Y)�=�VEjm6i�|	H{���I���]�)������:Fw/A�ƹ�Wa��S�F�w�p�+&���t��If�S�ƫ_m��G����T,����6��'��@z��x��Ф���0� �]���T���l��zIO�{�s�7����|��r���<$�r���Gc�����ɾ�F�@�,X�JD;�H)!+K������.�F�,N�o�]G2̮?��e���]��-�07�c�����(�a?����M_CG���Y�F�3x��1P"���ȸA��J����{��HkX���aJ2e�q��׫�E�W��(%�C���u�b:�qf?��|ajUu���@
Һx�*%�eT�����k;8�
�$�M�U\�,�_�K�^��p*~A\��#2��/���M�N3d�xK��#	�P���z0v#��}��EC��{�s�� ��|h�?��V�-���0i0�a�.�|�~�٠7
,?ɦ�}���J�2�2م"e��DYXr��R��e�>1����|N����� 
�=�6O8:J��C���h�ímoKh�
A�F�J�T2��c���w����c�J�f�%��;�6i����ڳ^����ۛ�\2�EP���h_�����6���/zo����\����^<��/2�_�1�-��j��b���A�����^q��vr-��hs������+OfW��b~g�໽B�z�)���,3�yrY��Rz�]P��r��bx���h�4'�ӇF��{�{Td�6���ݐ��Bܒ��4��ܸ���������M���0"=+f��#Ű�9p�?���G�:����a]����p��p����ɴ`y���t��e՟��h0El�Ѩ�AC�+K�pܲQ���
��d��!���zeP
Y��GS��@����bTF��p�I\i:�/�5A���٪͖[�}<�C�����Eou��݉>w��!/��Ԕ+�o�`A� {�nA����.�4:��� �{.�u)�>�Nhݤ?����	l%˱���=�Ά׍B�n�.��1��oղ���#x���(�,8�w�C8r��^�<�[th��
v׽���4�M�+�C�VK�ԫ�m��4���4:	!e��Y[� ���%%��yZ)_O�@�I?��-�;��Z���zE�ǸZ�<=EHĒr=R��K� ���R�Vw8�V����q`p���԰6��R�X�؃YOH�Gt��b��N<CC�V����2���>����ۺUk��R8;�Ӱ��-r<И�Kic��D'��P����ƉC�E̡ R���42p��#�Fa���}A3K��	��a�!s��*�b�->��һt�
�L����r�Н�T���-S~��3�B��\��v�.�_^�eb�Zc�޻���'`Oaqc!�y���h'Fn����J%Ġ~ 䮞<;�=pNh��%�xo�2��n��Mq,���X������o�H�R����]�G`���d~�K$v�#��;�����н���T��.Oqq���0a~;kԡg͗�y(e�p$Lg�ی��T<�
� k�w�Èg_�/�qo�����ڏ����Qiie�j����xu�F�c?�����L��E��ev�0r,��k�[ 3��5$��iȭ�3j]r!*�RX�ws�m����Y������وO1H*��g��50��`���!a��VnY��2A��n�2
�n	����u�9���u�E�ࡦ����?|=�!^2Lߑ�Ȣ���Y�(��/o]��.��Y���b��5=���ŗU?91F�/��<LTy[c殉��*x�ʲi#?�~�Q�X�nI�it��~oօ��?�Fa��iƛ������lU�79�l��w��G�T!0K��e�Gw[�  a�[���x�P� +h�r���j�nخ�R+��Q��v����h����M�q��$H�%֗Iqi~nE�"@'�cV>�Y4�#�*;/oڍ�$�f'bQ���x����r~ȳS�h�g����D�!�c']��_ÙoMrn�[x�6JN����U�[&�>)�wA�Tz���Q2��NP��|��7�L�]ƈgR��?�FM���湴�:+����:Je�'��<���>�f6� 0f=-Nt��^��xU�9=���uԴ���:����wH��Ҁ}JH�˰�ad�>x�T�w+�bm�>�̾�m�LU�Ud	@��	�U���	��^z�Q�ˢ���=�";���a�����䐖���\-��jQTG"�{���f�Hĕ�4���m��w�n�F�=B�d���0t�N%�)���#��~�cnC�,��=������%���-�F�J�a]*����A�Z���F���
��w)�
�zW�:�
ښ?L肉WO��'Ӎgk���x��)w,௞,q��n���s����WK2{�,��I~��SZ�i�) �9�^��� S�V8-<���O�����G'���?_揿Tj���u��BfF�:t(N.��y4 ��2u����]{q�ӌ^»*l/-q������.�8E�����ɖ����0��W�@�,���U��|�xA"��T�8/���I.hN�{M�1���	4L ܸ��F�Ra��%��>�6��P)��x���_�m8U����?i]��{��0�9I��`S��p�{��k�b���3������3�mk�2�*D�8Y>�����mAU���6�j�=|▘�� 5�������;�&⩹����Y���u��HdU+P�Z�27
��0�WO�<q	D4��w��$
hx>����7<M_�,���z�L�YP�A��D���=5>�d�NR�^P�_��:Kb��h��:@��DZ0zS�⃾<A����o�r��*�Z=����q1s���P�}�j#��Dn<H��Ji�a*n�D_�5��5:١X���@�;�Y�r���<�[Ǭ#����I����6��(�Ù�CV��]D�s����`B~�U��&o��@��Ѯh5�/�i�Z�CߒёU��[h3F�z�)��k��¶pN�)&�083B���|��A�11A&i���
�]Bv���zdi ��,d��$[tƶ�7���SxA�ʭ�%3H���j~#�؀}�~Q]d��_0ѥ�Ӎ-��^e�I��?*yt�;��(-JU��6$��2�A�A�S��s�wtc���|��	 ������mv�]�6��OVcњ�OO3��D�U�,]��"�1��[�G+�C���XOZ��s[�v&�{�"���<���OI�)�|��26E�������R�僥�3��P�>y29#&ԱN*rL�&�ߦ\��ӗ��<O�&�ߺ6���F�ū�&����ў�/� ��Q
=w1��y��3�tD�*�Q���0���z/#i*jM��Jʷo0�O-u6��MK�&�	�O�n�*f��誑4E�D��s���!���j�^��K�\jU�;� K�->b�k� >^䪦Ҡ�Ώ�dw���NěE�/,c��X��2#T͎rCO�ju������P;	C-(���cz���>\ \T}��Ȟ��
��!�Xn�Bz�9==U��+�"�)�.��B�mɷ���+)S��W%���ݹX�����Iy�%[iv7���C��'G�5q)"2��-Q���j��4I�ܼSJBy����G�q�I�܃�o{���}� J��j�&'���MӶ$�Š�]ù�o䔉C�C}w��w���G�YT���-���&�&�v��"�!���t|�`���feFt��5VW��'B��l
)O�,�J�Ij����Iu�S�No�8�	����Q�R_?���1CwK� `��iOlxTs'X�ANx�a�2����?�T��Y��wZ<�
E�N�|j���B%����ݓ�L�պ�?m1b1[�� ����c��r�O��|p�RV���.E3Af�?ݔE����S���a;��'bk>=���"��ֽ����M�AK���Z�7&�o��p]"���T�3ϛ���w�c�6�V��-���]UM����O���

����t`6��h%	�����c���j�^�Q��L`Z'�~΃ȷZd��q�G�����I\r/���f���@K�i�w�
���cqe�Y�l@L.�:�o�H��[�5���3</Ї�UE㒅���:�ԡ��:|�>���'�<5wM���
7�w.f�C���F��m��{�W�w��s�u���=��0$X��S�!�as�fF��t&�[B�P���n�1]s�T���:�$b�8��L�]Z�xl�@V���>��Z.k���Z�>xY%�`�y9�9�ܙ���YY�`%�4���E�¿Jqƛ����P��i�Ư���5�σ�ף�WK�&h�r��s�#_��s���~���Z��5Uq;������sI�\��;���ʺp����{ �J-�O[������Ώi̧���CI�![�	�������J���\;��k�9m�9���C�w�ym<�±pk���?�$��ƜK%��"
�t A?U�'Ņ���7&��cl��
j���Uև��}[�a������Yz0�UX��������
���kv���#m��/G'G��,��O�d�)WS4#=�$(C������M�@�ZE$�A�ԍ���D��#75� ��tk��U��;�����9 �n���L�_�-�I�2MMF�v/��H+�Q���A�w�_b�Cg۝zU��7Ϭ���Nr'B�,0��M��_!(����T�;?��4���5��Pr0
F�S���9�pG&�K��A���ޯg!���4��(�/��S�����6 v���]��7�Ѽ�[K�Z�N���%u	��U��v�4L��)ۡEȥ��ZB�Li� �����퇀&�K���UL)�[ ϧ��P~���7G�?S�ܯ�@����p�{V	<�>B� �\��Q�ޞ���P?���;-�dHJ^�6��Zd��xe��n	b��Hy�n��D䑾yE}t@���hW���O���!�g�!1N$��H�eO�DS�4B���\�E�6��a��f#	����]W� N�K�������Өm��F�ٷ�"[L�5������g���F��*��OUϻ;X����G���
�~��h�	},��/CĶcǈ�;��2p��>���ֺ�T����Z���q5}Z���L������y�ES�-xzR�9V!9���2����}��:��dW-������\9kX_1� b�����}$���)��h-�^UJ������[�e�v�_c/+Q����\�SK�u0T  +X�cZE1O���u~�ln��9[�pDK�#UU�G3�v�H���j~h�{��g�g��-��w+�똗���Z��������O2���ϽˮV�!V�� ʚ�����l�5h�V�"����_��cµ[r㑃��G#,�+'�Bd�[T��k��M�o�2d:��Bx��x��D�K�%��VhWSFb3kzMZ���,�6d�)D}�/�/���z<��-&��f�(͚�zG3Hvj�tÔ��M���$���WA啁WXuI�ni�F��c&i����\N���"2uÇ�w����Ʃɟ�����3m���O�i��������>z�ҹxWd#�}�Q�r���n\����f�ˍ�#�7�1Z��@a��s����_a�6\�'n��oAFK�(ʇ>����J��x�V|��f�̏��\ߊ�B�p���E�ظ����׶Ph�x�H�����:�4�qM"���k="�%E���*%�4�ޥ�ՉBj黝K���l�+x��p~M�a�3q�;��M�u��L����*���4��L3FQ���L: |�jm���e������M@��Q�LS�K~G�?3W��j���2�(�qL��p�X����e�Ż��Nt$ް)`�YU.#�o/4�k
O]�
���5���Ζ:StBm<���B�MbVQ7J�j��R}�f��3��l�� ��xV�xk|m�}?D�)��.O��O5;'	$i�h���̅?�zh3h����\p�����9�$>;<��,�/�o�	D�n����0�����[��# ���^�+��{�:�����Zg_�#��4����~R��^! 
Ҋ9�d���/Ei�v�C8F�ATly���/�ud@�w�Qg�������w8֞p��}O��)��o�sYW���ZjQ�������xz��/��
�^my>�W���l�R �~�l嶌1�	����v�vH�Mp��!CP��D�Ơ"8}} �%�j(	Σ�~��3�j��I��!�ަI����d�J8���sӶ�Nð"{ג�k�鳊�d����C�b��Fl���XNWd+��q~>{��*HL��-�>���7Ԝ��B��a�h{��n��!zP�=l�ek��7�n�J�:D�J0Rb�!h�|F{�w��,���b���r�����Jct [��r� ���~�V�d��Ǖ~�n��=�#U�H�ɽ�]�=���ۓ�fk�F��xz��BOdE��W����U�hP.4�>	`Sg���O� ^���Xcnj�a�Q:�Ff�OBSh5X�� }ym�y Rӿ�:d�6�)�u8]�k�/K�������UҢX���4%�P=QW��&��.m�uV���8rϳ�,_�?	4��u�CaP~�t�I�z�.oF#]5����?]ڪ�r7oi�S��7q`�a���jU�';���8>��Uw��̇�^FL�0[aa\2� M[�r�e��j�Jn����:g2E��� 7z$�2�U��s��L
� �z��b�	�����5�h�Ƃ{j-_i�`af �I����3���KH��B��o�����c�#�t��o��Ϥi��� 7I�Xt�t��ސW�hޠCl��ω`�@���+��ix�6+*�N6�Nl�����jB���Xn6~�Qj��	�%<����,r�j��xYX�CTY�g:U�wy����U�P����ߚ���6���9���U�O��o��>�pi+9z�74��@<P�'޳"$j\Nm�W�̡��^��Ɣ	]���ā�eol^���Xm������Kk�W���BhTD7��!voJk�xY[��ʾ���ŧM����}�%h}�bLN�!l�[r�*j;�_�?Y7�@ڥ�ZGkA����Py�Q�I9F�/~�4�w
�mg.BY�$�V�f�֜��֤'���m���ڪ�F�,D�9��F4��Ga��U
y�`��o@�ꩪ�'������$.����|�;;Y�˜H�YSH��,m��� V�h���S��ˣ�"��ƭ��p�ܰ@��o��;wb�b�9���,�[%�9�.'>ROӗ���16���"N�^��N��Q)oL�dx\m��f�4�{�k�gv�3� Zcހ�41jZA�"Ƀ��u�}Tf�B%:���vN�xݪs|A�:�6`�	gHx�q�iH)\���cċ�+;$<o4' ��2-5�h�n��{���7?o�35:��Α��8[� & ��C�DiRzC��t�&�����2����P"���bua�*��=@�Zo]"�zR�,S��h��hU(|��i���K�"�� �])jݚk��y�ݺpZ=�@��RKZ��[�������Ⱏ�j�����?�]}�t�;�]�cj�6c/��{�w4�&04�2�~P��#\�o��~���s�L9�����5�� ��b�c�)78F��g����������~HH�+E �}�R@O�����('�	�@�q83���VH愈e�?PU^����p� ��;Kxk�J��$o��[}M(3��-iT!7��:n0����������O����7�Q*�T����Hd6i\����S�.v�^_��<hŰ�9j/���i�Au����Ǭ�*��N�M�oz_zeb����D��M-���j�����в8k��5��.c�3��̋e�8rK4����6�>6?w"d��qWUjr�U��F�&�x�KN�N�_��]�υ����A@M���ȱ������pw{�?���F<�<'���b��.Z�a�2�p��DLIJi�It����}���r�x�Р/���
;C�})-�L�m0�(Ƃqr��	��NH�^��'{v1-p�ב][H:Fp�MY�[N�Q�p8{��n2 �+�`����p��A٦2w��O!u��;�����b��LO�R��;�hh�Xذ˫�P���	*��ў8�6z�� W��w&��y��O�f��d��Kw�G�w6���*����E��X@�.6R�}��pv��L�ч���,.־�S�=%�F]@���5���_@A����׽�{(&���f�5P�$G+����i�F�C��A��$!�$���#=��e����n�ј�L?6`��XlwIB=N�G���#�o����c���f��ꎕ�Y���F��A"��$.W5R��-5R������'�w�+O!Q_�6�>c���Kۋ�������?�m�wu�w�t�'ښв��A-�<���L���sg��.ۍ�laD
��̎|]����L�J����,ums*�t���3t�Wg��5�r�c�	ط�g�=LgԠ��z�8;�A��M��K�X�Ct6d���@@�%�'�)a�Kl8~<��n�䞲}��ΰ���� 
�:��&(w���D������@�g��?A���`�������g��ö�۫0=l�-¦8Ms5�3�^Ǌa]�鮠�B8���ؗ!(���13�p�v�z�U�H7��Xփ����l�xh�͝���
r\�O�ĵ�ߩ@�>�Z%�����"���ߑ����+O�˄Σ��������-��5VA�ťD��b7ԹY���a�����(ɷ>٩���F��t���R
��LxԖ��b(5x��c��C�lR�����*eS�Sx������D#d���|5v��g0^R$�+��1/��<�i��q��&43@��3f?�Ӝ�L�D]�RЄF}rf��V��<c��xN�7��_�i.�͉��2I+��;�w��k��׬e���s����b��J;�x69#?zk?��.2gMԼ��E�Rзq�[�۔�h�މ�D��MPt*���o�gs\�E"O^�4���s%eO��� �m���#%�o�a���v�y�0�>�[\T[�;�ˏ?���VBa�aU�7�H�㧆_1��:'+7��7\j��7aa�B��~oAN���#a���K.?���>�i�ڝ"mu���R'�*���.�j�������=rS��8 Kp�2���Ji��_ِ���(�����	����5a�Hul�FT���r6�@T��Þ|�M5���K ���ɔD��B���6u􄭪2��I��^����[�X��ݘy�q'�ד~���!��	c
H�������X�!������w�<�w�)%�D�5J0O�aM\��ƛ�����2v��� ���1�;���|��.�X�>AW772I4*��/jr�%R�{���~ L�qd�YWe��� ؼI7��C�U��GD.:?%>���}����b�Z=Մ�"D�,7=V�kN��`'�i�ņ��r����>��rv?c!]{��*f�$�Y�<js� �r���������0P��;����Xf��K���B~�7+���-4�ט��6Ye�)GI�,h� pPO�sc#��*.4ǒ�}#�����N��;
�o�g8+>0)�T�I&C��?iY;8�7�R�z����kw,7��t�MW�'%`S=�j掅і_[�6�!8pWT�-I�1S9��JJ	��|��Ty�������`�Wҭ��=Lna!~�sܰ]���m�G_n����0����sA��U͘Ըp1V������p>�d�4\Mn
�!*��Ջj��3�hTc7X^R<v%Wb�*]������ESkD2������xo/�_�pn�>��h�Ĥ���D�0�	�~ď�$�+���816*�X�dx�����~�8\%YÇ|�_����NrN�w�
�&0�HU��q����Y+:���#��Ж�������"�Y�:Ⱥ��ɩ�3�/\�d~L��n�LQה�@�k�y�N��{�ߩ7`2��q7:ߵ�t].s�]���Y|���	l��"~mQ()j������h��,���خa��G���2<�&��?:�GO�����+1 �x��t�@fI��nF
����n��gBԵ�B���χ�sٌ��4����y>�G���5ᅉ���H�9V��ƖJ4
0�v�
�f>	�����Q��!@���1x2l��_��}�����-2gO���x��E-��A	���-z�X
���]�Fē+�BW[�Б��l�!�^F}�SP���|����-�v�V��+�._`�q,|��+��9����y2��\�P����#�v�O�-��rfo�2����ֈ�|��b`�KϽ�]����ػ?,˰Z�=�M���bAf�ZQ.� �9g7��u��Q�+Xκ����b[I� g�q=؏�����E+.ެ�69WB֠��"����mq�9K�ȃ��7Xx��/��޴仠�9[C��E�E��OYL�&c��B�Q
��K�
��іɼ���&�Eգ����3@�Ĳp�}4@Y�䇂A�ؤ]s��d�.yH�I~l�M��c1 r�z��h����֣� #�"<Ҡn��A�TT+�z�߳��,����M�?S.+��ʔ^�ʭb�,L�-9��Ɇr�a�u,?�4�[������tF�/�m�T*�5�к�v���V�b����b �=YT%m��-��갋�Sob��'����E�,D}�r`��c<��9Ц1�����6��?1�{�*�Z c�o	��������T�砄���"���W���Z����%��B�uw�]Ӟ�@�96��K���k�eZ$N^�ؓӡVo#6�m��+�^�G��6�Z��O�!`�ނ��ZX�3>"��̄��xy&ݩ-��%���ZE�0!X'%�G+T�H�� �"������O)i�6G#b�<�t'��~KԪr�[{Lڻ#��"0l&۷d-��=������<·�qV�M�h�6��O���ڍu<[���N����>{3���5?"���x�">Xpږ�Ft��9e"^O��\��;3�Rf_� ���6.(��
s����5��֢�},�jiՈ�i�k���t>ƽ45��a/��S��t^����'�н:�H$�A֓��5��

�Xr�FZO�+*x�R�%�L� K��Px��(bm���F��y'�# 6�4kX��)�Q�����E����R���l��@���)�hlf�6C���Qfd��ϲ��G�"��b7	��w�����2�ޠx��
�� ��2�995�1�k!
G�{2��(}�:��i2��rV�{~��t۰��~O,Qλ�6^�ފru䴀Sl��=�_Dϩ�²mI<�#�f�l�����萂���� �`v�0���V7��U`ApP�>Ѹgl���MLq+6���I����]|�2��ݦ��D`��:��=2��b��2h��V	���Ѡz��qV��"�C�&����R�?.u>,�D�A��p^0˾;&T����EOBL���=f�6�ύ�B�T���`Q���E~h02}� [���)��֗����<|^R<�������D�W"T1����3����b�D��]y}ݷ�y����a�J��#jA� j�*q���a")�Yd�7H�"Q�%q�,�¡���c6���&#Q疏)6�ց��Rf�K����,�#�F�{��( ���VBo���SXYphr+*b���8!�*�=k��S�&�*X3����fF��a�f�}���
Ä?~�8�=-��*e�A���� �#9���Ov�g� yV�M-�g�fOg ��<=ΰZV�Ɉ���r�����ı��FG`�$^������Z;cmڧ��IT���p�ҁЇirH%b�:��{5��o ��業�I�7��_�w>�~�8%��1F��6��?�h���	����ম¤ts�=�5���<%��M%4����!h�-!�X3����w�<;yp
�����G4Hj
�~)R3o.��}>�U����t�3�U7s7�;>(h��d��|����i��_r0a�02�[y+# �\� S�����4;�`�K 5�R�g��#���l� +.=�k�#�p�%� �B]%�A����f�	�Nx��P7-R��2�STO��=��q��C��Mǘ]F ��{i�=Y�K���/�I^��o۪�q[F�V���d����b��ŭ��V�nZN:p�S���������_��P��Ҳ�4tpm�W(	��oY� {eE.L��}&�œ��������uO�i}��I������"Sg$h��$;X/�� �J���2 i]�U�.�� �)!��4�-N_"����=��@��	ϊD��A���e��ĺ���:�^a�FӾh�2�s���Z��Y�l��.��M�!�b��5��g��e��+^���ܭ��>l~�:���	�vs^�s'
�2���`�TZ#�T�:n����	�!�;��p^.���F]-d)�E�n. �F���G9i���S8՗ǳ�g!"�u_��X��7�_�ER���-9)�f����>�B�H��V�jU����gڶ�Z�-����z��F�c�fD2s����e";��2���. 0�4˃6�J�S��m�Oŵ��%���VI_�Ջv+��\N��,}!���>UɺC|���i���i�2�B]:j)���8@j�J˥m��&>B�[l5���t�	�c��?��p�_��}�%sb�H��xoBCW���ܧ��E���C�m���F�����P$b���)\�e��L�Hl�5��֗�������M�����F�)j���d���7|uXDM�&K���ն늓��Α�&:Z�5�5y���Ѝ���f����H&z˺g��^��wku�@�T�	������j��6p!���"d���ﾥ�9�=m[��^=D��Ν���h�!��Fg`���^��oJ�d�I~����s�X�hŐI|U�cD�<�h{>A�})�ʙM�(M���}-�+�J
	>\]��O�������D�=ڔ�UK%u���a�,��v�r-�a��:-x ���Pз)X�u�V����tfY+/>����喇��겞�\�9�蘉���N=�pA���\�9��Y���G�+��w�� C9�dym�0TӁoI6����)�������l �1'�~��}��%�'�m�ܨ�X�%��oI0�O}�4%�sP�T0;����\#����	�i}뽕����O�m�Q
ȸ�D}�|d�^�:K-��b
��8n6�����5���)��z�7Q�Z
���O]D�e2�v���%L��\T}� �]0��AC1,�m�2dz�L�W��H]�<Š��g���0d��ɇ��'k�:�C"RA���F�+�yԱ8��<���{8\��N��}����O썼��j��8g��%�����=F��AO��t�bh53Ff������N�IW�L�����.�L�q3�h�	ӈZ��ILO��#��I��nU�ge2l#<.��� ~�J��?�ޮ��H�{>T,�ruŃs���R��^
�~R�g�iߵ�ɥ)�&$��.@���[�KШq�T���ZMj��8��Is��Θ��g ���㝖�W�N���
x�l�AW(���ٿ��\�RZO[���o�XT ۰�^��o��KiLϝE&x�f%h�9�)�Yk���R(=�RU�bճÛDȝW�T��b+�阕/Ǟf(Oy���~�uS]�NU���pd�ü�$�J+�&YFq�(��dqR-�+ ���9U����(uJ�%(a^%�:�SK"#�~7@�h�g�����Dd�hإ�<2��M�� }Î��A-����7*�=�!����O�f���9U�]�OK��ly9U����k�
�ȫ��;�b�Lף�!��%z��gu�ծ��u����'�o5D�DWº�E��X�y<�b˵�T�� ��$���B�������$��R�VI���+�鼾��gZ{djb^y��h�P3�	�ʠj'��n��Vh�E����,���"�H�Wod�'5 �kZ�2��q?�Ǖ^�$
�
`���-ȁ}�`��F��*<��&q�X�r7eYE���v� - {�r�;o�%��Q*|7L����K��rX̓��9d>�&�~k;+��H!������)[�'��Z)���vvޔ�"�͚�MI��:d"̺6�Wp�b��_b#�X�؝vA����4���	�n��2�I"[���]�����5˜X�{��J@6�˧p	)������|L�.z.�ܘ��ͬ-z��j�%��ywR�k�Z���"�s"�׭���K{��Ǌ���[
�޳'�X���k}�|�޿O�(Z�^�td��d��\}=�[#�_�U�pϋ�-M+~���O������k�éw�8>��u���$�_׾�	^ّ����L{}mw���ު�JŠ��S��fC=�|Խ]���Q��վ��k;u�0D-Km��>�[��ܡ%��&�������XQ1�q�zPIo����EO���8�5�Į}䜺+ e� :J�l�.+àh�e��/�g-˃<�*�s��&�+�s����P����?,Й܆�EIs_�������rU�rI@�׈��,ZI��~�v�]wu�R9�J%����Ky}� ���i����՝�,<Q(hf���.�.V��]]+5m����UK��L�c)��3��l����z�U�C�Ti��~�j���DD��܉�dv�,��O&��`�wgi͘��x[E�6c��=�lT���kӨ���G��ѳ[���'�>�^�F�ޢ2=���N\�#KYӒ��)����b!D��g�j��w�e�P�M��H�R�g� _
������\r٩�͗'s���8�jA��90_���ש�502���� �I�{�=�����G�fY�_��B��7��B&*A41���d�WCe��Nϛ�0�V�S��~�o��B$��t5��iU���$qb�����.�.,�}C�#L�����YxK�ν�-��r�XX������پk�Ǳ�8(����\�7UNcZ�R�4�6�Q4�CrG��|}
S�iX��M	c�[2�fJ���=.�VP-2ͱ�-���k��v�"��4��r(b�~1����NHC"��<�#��N	Q���j.�#���6,�w_�?[ �4]�5�|Y��ℎ������J�����5���X�Q<O3��W�7
1�Sa�==�ْ^�{_�;hv9�2�| �H6�)ĭ��x=��P0�d�ا�|s%:�+�K��]�0�Y��8��tJ�Sh6H�,<9�u�Āj�	 ���4[��#�b0_w�l��� _��|�����a�w���V�����]'� {K�[a}�9(�
M'l���1��*^g��~�A�W����p�ꝋ��$h��o ���+>f��l�dH�0���N�ъ5"�jp��{DPr��/��p+�J��o;o�K=��� �@KY��5*�wvX��9���h�[/k��]( \�^�E� 7��h<^�m�["?���7��z�1ɳ�mc%�[Ɔ��Ś1���BoKi��rUi��E�w�@����S�����.1�kf�B�Z�;K�����B蓏�4�G��"RK϶}|zY��S����K��+3OUMXU��k��7/�J��5>�_��d9�j��jzQN�Gы��E�1�]$eݹ8|Kƚ������$3e�.�_\?�+W���`o�?���G :��ɟ˺�~�?�d0Oi�ۧcV_P��pl"*�b�U���4��W��@���l�
���.���+�Ⱦ���w)�T�%���:���<��s "ͤͻ��i"�f���`��W*ͥ���:9�(��w�`�R�&]�����k r���F���7ל O�i?�`7�2k8��K�� 5�_x�|4.>yl�����<��������fWՈ���L��+�cH�3���͊y�J���[T�	պO���곽�S��l�2��{����ܾ��+�j	��G��-x�qj:�gq+=��W��'Fk��NԹ]յ�?��:"�������ǀ\�9��[�b5k�R<�D߯H��.�W��ٵ�B \܄W�����#<����i��ӎ�#�5M3F�ˍu��@����>h1Е��s�_ Nfʬ��Ĝ�}�Bm����=��26J@�n���|4<��p��/����I7�(����;5��F#�H+�+�$����"K� 6�Sr����W�b"^���9u"���J"�k1ǀ�k�f�K���>E���X��4���+`� @J}��b�[�xJď�����8a}�O�u�m��Y���#P�G��ѥxYD�yM�K��3�f���6j�g��_�=<\1Jl�8D*�*�_��J3�M���B��|�]�w�!+�O��g�Úh��J�ͽX�����������_B� �鼰��l��Hh
�S��f�,EC��bZ�m��3��z����`�<k%�M������L̝:�o�u�4%�UXA���t���Y�&��D8\q��y"���O���@:�p��CE�`/�۔�L
[K�S�^9hB�HX81ˇ�-�m''�� �/ U��#,u�>��sA,w��6j��H�<�)��߷;Ll�k�u�\�C�b��^]y$l��}eY��.��7O�~S�\�޹�3�|ާ�	�PZ�,�h�=P���0���v{9k,�����23������7u���m��S�1��z������y�!�����ź��;c=�We����Ӕ뫑�7���|�8[{��0��ۏ�4��[�j��Y��DH�>��]��;�2=���A���B���Ѭ�7��q���!��/����~�~8��$���Kˊ<��v-
#������н����Dl�&�Y΁�x̔���p��j�-c ��r��^�{3�ņB-�hʍ�$�A�n�ue��D?V�q'��+Wo0�۝����O?O1|�x���Wnc��En�-�R�%D����;�7���	��w=
ے��g�O�HϿ�jEw+���w�]�.��m^Zu2\ρ�O��e��&���xS��(����o y2:������W}��X��#BE~�9��/����P�k���C��<d�de�B"�d,0�E*bvg�v�\�1U�/���/d�u�����ٲN�l���ޭ~9{6�fM�K�1�<:	bT |�e���m����n�L}��0#qձ�$�溯�ҭ8H�Wz7�mv+�������L�%�2��Z�����x���Aڿj�6�l][׈N.Pkz��r�L�G-��y���1Wi��f,�NM<�]���I��a��Mg
��/�_f��S�7��8�;����.���C��U�t�C;�m�O��q	�: v��9�7qj�����I���g��^$�琭�� ���T Ӷ�QX�j��>���}�G��~M>o���^��� �N�����?ѿ٧��'��C���\�a���m�W'�/���w�`7�Y��>�.��7�ӓ��B�#��W���>3�"���u��}�_Vsk�a�5N���<�{a1i�B����
��ݳh��H��}5��Z,8�V}46�V�A�5z}m�*���@���x�"+W��j�X�Ⱦ$W='�L�'t��!�G�-��.#~��L�K�>��
o�@����4�b��������@K�=?��Z���c�I�I1,eA̉C��r=���x@h�3�!����rK�G��1kKD#�C~�;��+Oy�)3-�&��@�/qIi����TM�G˒7-Ǧ^�Tۣ��T�"��`�6���J���?1�o��p�Y�wE��TUP��q��|Y������&�'/����F��n��4�';غ��_g-��Z�|u���BI-c�����Qn� 9�S����:�o?p+j�1������7&�{}�	S���=��˨
�GA#���5ʮ'���k�e�ɍ�Bw T��m���yCto���Yܾ"m�g��C	3�-d0U�����L�{"�B�u����q����}�R�GX�]�"���yTD��t_�B����spu�E04k�Fv�=�_�T�&��h���~cB��(
J��O�Y�����{3�'W��FW�0X)����ߛ�<W��܃g�(��[�`�_���{���0NB�ì���,�2�Z
���7������ ���y�hk�z�/\b1q�%{�{�A�`��Ђy����M���.�YC���"��q�b�b�vׇ9x����0�=�<��HE	��|���Jݥ�����Ļh�F��)!pv�d!A���¾��>!�8���Hd�;o����Q����*��ױkIJ#{���_�5�,`��E5�fk�ͺ� _MT�c�6�Eʴ�dƕ�������%�o
�e𑻑�{��K�ʃ����{�}���"�hxܩ���J����u�J����� ��d�{�|a��[�\�pU�E��@��c�z�,�6�c���h�D�6����ڟƝ��9��	�9���@/oyk����,�B��c��@sQ�EF���nˆF\�%�ϋ�Kd�Ƶ%�p���ȁ�{�D�?#�&Hc�T��e�A�����<k���Q}��NA?�Fh��_���@V*�?��˅m��>��\�Sv���JI�N�k��᫻��S�c�ɎhBd�:�����UYx(t���ì�T4ngUk��r��;<U�����"'�irt��@��ڀ%�wɒs"3P��DP�
�QZ%a�e�_u��e�-�'t��p��L�]��X��#)�c/�����!-mH�x*r�k$H_��*�o,E��l�c��г�"��=�,�����V-��ς�_#]dj�#c@f��#0T2"�;2��,
�Z�'�<C�@l�.�$U�������3���f�Fd%l���
;+�=�Ԣa��J/�ߞ�zK.�D�7.ᨈcK�Tc�	��V�29�H:u�)����w�{�;�RGϻJ�Ѻ�j���(zp�'����4|�Bȟԗ�y���*'`s����� F�Ԕ�E���|O>A܎U�k��uL�O�����ݔ�d�e~�t�e�Z׉�4�t,f��)��$P�*�U�@gC���"���.����9*��M)�ܮ.!��	"�S�'�ܕ�2ƓX��G6[�����|����D�&�T��.)�/r��)��vI��TT^$�L޸E���k��@;[����iw�����4�7d�M,Ro��1_W9S��H�>O[�|�M����%[�������Y��\���o��������xe��F�פO�cg^���H��@I����[,&�Ml��5I�=��rբ� �h��i�;M�9�ƐcrپW��&��q�{r_��	�7H�'�!S
J�P
��2S_t��#!(�?b�E��t]�����ፚ�Ӈ�ƁiB3���]����H>�o�X�4_��)����#H(��>�	������.w1aM*w���=�s�2Y, ?;:wU��RI�$�yG�M5#~�#�1r�������
�V�Z��H�����l���_�/�g^��/7�e�}�F�d�ى���N1�%)R�}ː�I,�8�X�K������;X1��2R=;-�#˝�@�'
pP�G]���..�y�=���H��O�''��lv/�燭E� ��y�p�R\�����1����'�Y>�tԉ_D��k�ݳ�"gT�]IH,}Z�;�ߕ�XE̻�X�掫{�_�ԝw��Z�Û��0��iKZ<���D���r��7:R��_`�{���G�դ}��=�΅Z�j�rkwĎ\�8�l@(Tߎ�O��-S*/�K~gy,,��`����I�M�ؔ�|R�v���fU�Z��.���A%� GI�|{<����*��&�B:h�`v��t}%����̹����۩AY��%q�R����1
p�b��u��#�e�H��M�zl�g�L�J��)�����
�*���25�0�o�?�#������P������A�8s�k�M�T�ͪɼ�x���^�0��N�`�@��� �ފ:
�8��X���J��ѡݽ���#nz�	��m��f̕O����y/�,{n����7���ʗ,8H�D-�SH�ۻ���ǀ?#T��%c  �ޓ�����s���|-�3�Px�4�2���;�~6
Ldj�Z�ی!�Uy,c ��Qǐ�oT�Hv��r��W�(l�!)Rc�]�O��W!%�M,�
�\#�i[�|�����"q�J��fԏl���&�/b%�T�h顀��j���fO��\��ӊ�=0g��3�m�����i��3/�b�&��`�4����L4}�wU����8�s���O�� e���	q�2�sk�d2��}�2��8T:���h%�/�����^i�1"VFB}���%�����Isz��s�~�ܛ2@(����!�4�EU��ʽ,)��d�}��wt;ke}�dc��_0.8>�!��t3}ڝb!RuO�����G���'�Y�ӊ$�x�J����%���9G �C��b�=d�b�"��"�뿿���h}d=cW��,��O���(|JS���B�Y�R���ul� CC]XK�-�!~�n���1�J�4y�'��H��F�#8�[���T��;�����V���]X�Յ����^�`�e�pԺ�E5�Ro^&����֯�Ӕ�!;q�e�=[���i:.����׽Bd�6�i���6�U�p�d��d�'{�#R~����߿֜��ͷ��m������x�1��<~Qɲd����r���~m�7Y�xK�u���N�C�9�����@����D��Y�F�ۋ�3٤76���4�����d{|1���x,����e�2Ue��b[�|,���t���J�sp_��Wjۄ�u6IψPp��=��#�7pa���,�f�P�a?il�rͣ��G�ɾ�(_����S�����W^(�=	áS��fnZv)m�\@����q��պ��lO���##X��}�vp��1��r��f�������tt���5\4�A^�}ͭ I��U1�u��6���92NV���:�s��v�!��d����U���<��6.%�[	��H�S��M6e�8�	���);�"�� ֎YO�ku�-�XG�J�]�`eQ����K��2sf�\�[E@�N�i��^-J�\�Iv��.���`+��%�_�Ym��km�Lo�%�7�#�����1嫑Pm6�o���;��+��ߢ���`5F��м��w��j��O���`ߧ)�> ������=^U�,N�z
)F��hrC�q@W�A�W�����у)gk�W��h�`��
����a��]�z�u3����������F�{�d�؇�&_b>:��W�z��g%�A
1��C����ڃ>a��}r������� �P���qt����t�%P��ۀ���I��{ �g�u��\�_���\@b}3��Խ�2��c�ğA�2� S��
�F��`��%kjUG�o8�}�͸�G��K�3��l~k�=䀽D����Z0�h�h�x|��������<&h����xr*���q4��m̹����^����.Z�B�ua�9Յ�"�-� m�5��,>�x�}#�]9O�0�G�:�lR���S�U59�k+���R�2�q0Y+��w~���,��9�(?K�HY�H��B�#���F�5�_:���Z�+�guO���gC��:ހ��Ź#��t�!�rރ�fh-q��u]�3s��+���X�Gp���y���.���O�P��'A��[\�Rj�aR��I'��PSc�m�\���]b�/�Y��œڿ�rtC><'���Y:9����%̟v7~�"�,FT��}���I��(�u�~[���h�D�g�M�*�s(}8aѰv �/viM_���<��Qߑ<��|3ۭ �D�7�݄�c��$��y��U{[��X�ݵ/d�5����u�� z曥�A"�s�����<aa�hd.j�g��?ق����[�GtV,_F��zOz�]�,�߭�ӭ�ʠ� P�2A�R�6�^O�km@��B��ZI�2tE�ݖu���ҿ�����J[(����{C���� %D�)�������x���� McG��}e�3���0ҝ���9�[���������!-"Z��v�SAM4�~��L�U��}�R�q����^HDE��.������ƺ�G{�h_�I>8Vi��R3w[��`]�nm��	��>�tiW�g��Ǉ;�I_U�)�w���cƘI�?�(gU�	H>��q�=�\]u4(n��ò}�O(=i�U>��TK�ƾ���_G^�|۸I8��I��[6j����z.p� �?�3B6*�<�׬eV�t �|��\`ƙ2�Z�����@��$��e���A&�{�TK�?J/w]E�cǿ��:����� #�v���E�Y���?��������|1��C�O�U,����f�����<�I�";��(]�߭������br�S$�����x��T�3���1�ҙ�}�Ȣ�!a�N���us��Z�V��r!�pm	]חj���}�DB�%�������v������F��^�?Cח��0�Q��]��9q�,��K�:����ri"'+�!�`���L�L��)��kt���#栲e��3��=��q�&�3��!�?�k)n��ٜ��?�O��6h^�-j�����7�k~W�\h��8K�!55ҦӜf� ѤӔ�3�n���xo�Gf�/A��xє$��i�5-]<�)�g-QL3h���Wm�Nt�6F��3����]q�)k-q�H�q���F86L@wȫ�V������PX@!�}��u�p� ���"�u��dD��sӣ5�l��^\d#L�f��-���D�y[w
F��͢E�����D����ؕj��.�q��/��D���ұ�0����5�Rg�Ź�ʥ�Lڪf���o���@Kh x��i�/W�E4 B=��tx�;a�8Ei��g�=txO0|ޖ����l�4<C<Q~l��Հ��.�<zr��!-��g�LLyGiq.�� �Z�&g`�<G �y�� {q���&��G��Q�Ykg���z�7�r�]vvȻ��U�J�[�#_��<,Kr�ّ�Ls�U~5���+�D�\�7���w�q���YE ���5���*�L7H��qӏNs����p~���:��"�>?_ڈ�L�}�42h��w����gv��Jh�" �A6�׸7G%��G��#C��	kwް�h���%�k�]���I��ڜ�;l��xD7r�:��'9>�(if����o���Lެ9�7iC]�rV�24�T_)���Z�K$�Sj�u*���քF��֚�J��\��<O�i噙~��3務KG�mi��� 4� <q�"�.f�Ѥ֥\�W+�	��V��_b�}�*�Q6B�����K~��xM�|�e�Q ���w�p��O���o��|@e�ԫ0K�u��=+���h�9_rY�9,�+f:��.k)��y0�e�d{�C�����Z�YiFke>� ��'m]�(���8���AW�N�Hn=����\C'��g�j�����َ����cw��~E0K���J�I*D]�sm�]H�hj��j6[�x��δ���C�uev��Ƥe�s�%�,�n��c��>���#K�c�iL��9S �|��������*|�%͆��9�t7=,GA����8|��6I�Y�xRŜH�U>m�AT냺Qв?&F��T��WvL�*ꇱ�ܷG[��Y�Ή���Ѳ4B5\�r��꺽�]�,�T괆692�q��U^�wg���7!0�-��$�J�@�6��d ������&�̣;'���S�q�$|;��m뉜B�=)�HY
�5���o��>���d�~
��O�_>u`dx�TR�V�u�� ����݁�a-k��f{���m}՜p�4e�k9����N_8CG��mF��Ɉ��qЁ] H2<�}g�O[i�������t���FU���	��t�X�~��)���+!6i�7D��V�Â!M{`�Y�FY&o>��y��g>�����2�7�� e�1!�r�,�K�gi��d/�޾ w+>�T���ש�P{��ȷ�5�:���"�N�~Z�	�O��ϧ���8��{i9+��B��Хk;� �G �Ͱuh�3
P�G�K��P�#�\l���i��p|����ӆ�Ʈ�36 ��R!�n<6�X�E=�k
�'-�4��׀;�;r7���U��j{K; z�E�Tju�q����2HHUm�(r�@-�r�P`�K�%uU����� ��j�L�{���~i�v���u�b0߰�A�SV��/�����ӟt�E�4$�����O�a�dǗ�x��q]Ҁ��5����*N=���c67).��?#��ꅍm�Ŝ��{��6A9rڿ8)��xN����Z3~18�U�+�OSD�z�7�/��M�\�{�۞�@D!���0��� e�l�y��]���*v�T�	M��O_+�9����̋8�f c�ҫPHۆ�3�>*��Z�?PX-��ؐ��T�g��4���qϩ�Z�Ec����G�J��� �bgK�Dn(��j���ʻ��Ϟ
��dX���9�i�w���}���=�/�$���/��2�%�v��׋���tS;=��y�W�&����J#�"�8q��8y��U�=5>��DL羽��cZU-����X��1솚�`���^8���IQ�./X��K�{�HlFM;;��}�:�_2�i��w��@�C�d며�8���:�lI6��S�i�@����n�"Q6W�3��[�Jd2�kܛ�2�!��D��k�f����{^�`�G6�C�תS��¡~�1d4�%<ʁX��3��6����uH�cȪ���``Q��[-c�c{e�`>���nq�L�&+�X��A$����"�-��Z]ex�� ���,^~��D)#`��5�+Y�Iu�bɼ�,m�� ��ז=�	�9M]0櫞VED�����
l���g��(I�@dw��b'�Z�)Ҥw��Wy�[Je3����c��0����B��؎���}#
��� d��_ik�2HG�<
�rml����-�D�8�n�Wh�)Yq��ߏ�&�ٗ����nS���>��B<�VƂ�Ռ��<s/�s;�fc�Yv�3hyH�1�Ԥ�%�ɣ婁p5���5��	���#Ú��|��h"�M<��Ѱ�;#Vƽ�^"|MT���J��O���ɁJ�j�.+����X������ت��#�d���ZK��t��*qJ��[.�X�hԤ0�N"v;��+�e�l2RJ��57�Ym�=R矞��`�Ҷ�(���?r](����ubN��|��׋;��t^�ۃ���%���V����W��U���ϩm�.�4�m�z4���_�n{4�R	S���u��_i+�o�n�OŚ�$ʹ˩��M����y��3a�=����;�vU?额ta�%��UMd�U�6����L`�>��0�!]��}�������:�6Vy��p���Mh�`��#�n.`� ��s>Ȫot��Kʙq�<�X�	�����!�t+t�̸�52,Y۬�m:)(���5	[L�S@T��FjZ�U����*bΑ:�I�7����7(U�[) F�:�E.~n��)�ih�T�jk�K���_�m%F3k�'%o�w����I�|ٗ+��GS�H�E��Q���ڋ����Y���#M�-�!�FK��B�{�'�����\C ¡`�e��j�COO�-?��6���AO|�����U ���s�YRY�	�Z��Pw�܇����Y�<(4�CW�r�f�m.h����I��o�6O>����>^��'����T��v��?�Q9x�%�\N��o�UP��p���d,�TxW�aa]"U�]��_a�H��L9���J@�������<�KXoJ*��H�b�����1�6�.Jd���
rs�i,���E�>Y��˿<�F�u�l)|@(���=������,>�� `&��)?��z!.���,����v�+O�9�Aȯ4�:q����/U҅�#,�;��@g�/1��Z����˯/y����B}%~p�_*!�d��WD��Px<���٣k:�e:��s�[ەEC��XԦY���	���4���$���[w9N�p�g� �(�}GZ~Y��n47jh�v���vc'1KbG]i���/53�%BT��M�Y�Z�,��Wr�i7m!�W�
�w�8��2ݽJ$��h�4Г�X�M����|P�Qx˷qGD�"(F�*�Go����&/f;l�و:�8�U1/��Q��׫�/t�Ѯc�*pʻJ�U��w��1a�G­��M���L��^���},�&�P���>ڔ����W�G�{��[���_���xK����$�gf_�[�J�)�a{P�B����bzV�`~�z��5������w3��Z)`�� ��vD�x��!@^���Mg�rR,F��j��q$lOh�����#�L'([!u�z�w<� ���k'"dt��:��t���U+���h�p�����RTgLXs��4�zǪM��Nd6c�K� %#�'���FDLC�xFވМJ�S�ä�������H�R�LD��0#��;�B���ԠC!L�$P����o��/\�]ƾ�� ��q��V���Ӟ������rCT��V��;�G��W�f��9��ث6��4u2_����:��Y ]l�D������d��(�cy��<��S��=�?7=e4�wȁ�)� C�Q���h��5;�f�?�@`��jv�����hΰ��nT��������j��nԪ lb#P\��U�*=�Iҕ���j/&'c�.�^Q�_�������uQ��=��K�VY-po^]�T�,!v��6gG@�E�LЦWϱ�N )� �u��X[�Q,�3�H}a��e�@��������'�i}؟v��rl�Y�W�ȞF��fl�[� �n����-��C��'��E6#y�M��.<�^��ZB�ݨd���rG?����K�":�w�����3s�R�,b�������Bq�X-7�<Z��2�N���A߀N�IÚ�m#�9af$2]q���tS��YF~�d}�3����&���|�ϻ9��ݺ�1	J��9?41�[���I� ��՝�*�G�Փ ��t�S�~�/E�E������	%l\�#����>�-��G����胤�$�4��D��x��^5Z+�����?{t��w�����%��`�ӹ�3�U�[��($l�Ό��ع=	
ӥ�<<�a&[��^uL��K�"p��c
c4�H\��Q y7���N�����g���i���c���9B��1�j��6�<��/�$�o�����f�OC���c
������@�H�\E��T^�񳏀Tw֑�a����O�8�� �)u*Q b|/�@��@��<�oc�A�-jƐ��&#6�����У��os���o@j3e�m�����������-8�i,�UJI
A��;�� ��m���穓YP_�N{e�zW��6�7�	��S��0�v��t�=���������`��5��̈́��
(g�� ?4�BY��GWH�W
���,�U\|a��D1J��!�u���VO���c�����=�oH�|������j�(y�`��!ހn(F��I�k4��OtD�vSB�\�J-֙���t�r�K$��">��K��Ք�HM� "���]Ėe4�|�q7T�YT�(�Ņ6�4M}�H���v����/��OF;��m��7Pz�3~��t�*=�������5���M��3i,p����.�)�O�͚~�Nt4<�67��ۮ1,u�U*{��'�Z��3���g]c�^;'ysP�U(a�i���||7�T��Ͻ�i���'V/�o8`b6�q��\��
0 �o�x2�:頒Ό?pN��։
�O�P5��)B�f&�]���Z�-�����ҴH0��L���7�˼&�&Z�g�.�n�~�!jX�dr��E�z���s��鯾��n�g�>ݔjPm��Yҭ#��F�sHhJ|B�����;H��6�ǻ�
h+��v�M�`������I&N�LmFZ�#mW��UoS�J��3JQ���>r�k�i�eA(��Y<Jy���c��ٿ�e�ɩ�z�ʇzU�DG��ۆ�4~�oZ�VJr�p��%} ��<~�HoG6��k
×���0�	�w�_z�H�M���J��O��H�_NQ��w���<z�wV ��n@���e�h4��.�:�b�\n�P����״*�Uv�-(�j,Ԇ�y�BiMV"ϞD�
/F{��"�>n/(1w2�eJT��	n��`�n�2�<6qG�W�S9��'��(g�A�� #9J����j� �|=�C�G������Uh��Y���b�(�F9c��OgwP�x ��
U�D�,&6��
�uw`�KDg�����7�Y>*�ٽMo�k����Ѳ�n�F�8�K�~������,>�7'��L�`����9`)r>bVƂ�y���ЎL�$�3���-�a�����~���X�ťT�Dd�tƻL^����T�P]�_\�0�]�3����X�W9�IE��Gg�_�oF���[{����)�����ܰձݝܝ�A*�O�b��5�[�y�7�~�P�ڴ�?�0�����|����"��T˝MX�6>@V`+�XPq� !b����ؽz��J(Ӑe��c��9"���}�D=':e_q宄�%}���o�%=x�:n2��i<@�OI���%J�6�1HD #���eT�H$�΍���_��T�&����6;~�bd�'`�#1�H�C�_%y�����E&��v��I԰�\�&�T�7��u�[`�8)Z{C�V��6�/9O\(��qOr$#H���M��z��ny���[�m��uɧc��+hد4���W�&�N�v�ρ���(Q� aߝL��7��U����~�m�*rl��h�>2����[�R3瑧��c�-T27[���콝4��oD~Q�]���+�_��dm���1b6�h�b(��}�| $��$���0��O�{_u؉��"�(ZwY��y8�|��&�����މB�����BU�K=+�i�F�Ss�7�u��Ċ?�Ce�
��:�q فp��':jv]>����Bf��2��E�W�yd��&Tb2��IPҍ���ԇ*��6���"a��	Y��f��R�*�|���x=$xN��>	�&NG�F�k�M�H\_���d��q^Z�|ī3:VƋe��V㕦�GoӶ�G�=��0�'*%JhR���,��N΋��w(��;j�q�9Z����K��Bg`H���Z���%�/����Q�� Cw%�W%��Td�e�L�	�je������@��C��o W`Nd�B8��T�T���:�8K'��ɰ���o��=�Q�r�P���h�qր��}��� a�l�{}��pwT� ��gi����b�P� �����YǇ��/nS�+r�k9B�-�SH� ��/c���E��΁����E_�W>~|o��#!���f}O�z����Z��|���Wc>;}�����f~�_ã�!~�\����0�d+�~���M��_7����U!b
�Aim�N\K$r.*���$޿�+���n� B��?�E�VĹ?F��I{�z������h2.ʗ(�Vn��lV�H"q��%$#ɰZ͊i8�'���*�d��e�m��E�I�b<P�/��D���ʼ��U��b��WW�l>W��z�ű�.?�����2�=�M)g��������93�69%_�b�#���I0���GK�Z�ʗ�x�*gͳ����#�F�_'��	�ҙ�N����`T�<�,I��,��`&�V��+[��q�a_�t�w���I�e�u�����ɖ6�������׍ȓ����5P��w���	
��jMr��o�B��I�7nW�)�}gJos%�'����+sH@E���2I:t@��Qj�4T�u��b���H[j������AB� b0�,D������O���Y������q��!�Φr�)�Z+N�f��O���4&c4)�80��<����'I�kocV����p���
ŀ"�7���(>��8�P]	�ƺZĊ�k!��2h��Ǯd��h���:9� ��ЂP�Q�[8�8�a._r���6�����a%������vC�\s��Z��N�M�����h�"��˟��z�o*4���f�?k�I���2�'�cl�>5$u���9@�V)��#�rxT&���km�v�l#��"�F�ܐ�{� `W��
�hX�U�{��j�L��)�dV����6�pJ��8%Kh?���� �-��{�W��_��M���c�t��VX�\��G����9�ʢm����٘j"�rءm	f���z���B�;�8�����At7
�	����z.�4����IO��m׌����J��79"���t�b��$��yA����j+��K���Z%��k�XK��m��J�.�VVߏ��hހ��2���&F����Lg��N|6����R�	�>�������}���BQ�b��:QB�;|3c�G�����):�ъ��}���Br�_�g��\h
ʔܚ�=U_��{����^p��-�T�#�/ǭ��p�����d.E �/�1����Ĕ�Jvh��-�u��=����MY�@�pJ�7�Qy`{�+�s�.q�?�}P�S���z��7���m�2m+��������f��	���4��H��B�f7�rU	l��4�|�Y����iTr������`����R�F��U��������ll)z�Z ���s��n6�p��r�{H��7J���T�>=�m�M K#�R�P
���@x(eU����j�}Zv)/��.//
6V1M�k1ok:_�ѝ:]�c�b��v<>�%�?�A��D����N��Za��89e����������������Z���z���W�lT�H/4���.fn{����CD놩��F��g\�C�:�1��1�������#�,Z/��ٻ��%�&�[��(������>6�ER���4��K�����G,�,X����m��ƌPy��P.�d+�7��!��o8Yǜ�[:�"��@�L�Ƶ��"[Rj�Fe��Ѝ'��	�N������"�!j~�����xF0_��q���z�W��&��������7�C���O��;��)�8�b֔nu:y�9Gѭ�hb��)F��<Q)��h�T�{��.�����)�E������e�F~�����m�ݬs���RL���%���`@�V-qua��9���#����ǎ�����.�������7ն�De�����z�ǶJŵ�T=;�%r�n�KB`w�i�
�h�\%?yўb�E��cb|!�f���
Z�e1<�\V���P�l�^�;�T��=�P����Q��"Z�m�9L�-�H�2y���L�lU����ls�:P��|�藯[��i
5�2@�|�+���I8�п)��q���B��4�����8V�Zxz%ɞ�*������M�H���G�P�<��oMw�1�~_��MM���f�$:aJ���	�"w�c%�L��$'�����s,_��֙Z�Hխ4��v�-S_��dEg��[2��m@}���@� ��i�$Śv֭��׃=	E:�far;�.��(2��~���7!2�%�T�,�w��q}�����PJ 
yY�=�����-��~%��� �����7����y�zxR�����q���{^�zlA�fu�9�5�I��*R/%�?�A10�;��ܔӐl��&��l���lw5^\o�
��]��'�,#���A[�]/<r"B�D>��2�ӈ���Z^����P�j@�ӮD��[إh�˳Zc��Z���p	�Y�˧6��iX����Ͷ�"6J�a��p���$�W�!��{���4��CL�z��@�>f1�|)�mG���')���R�u�!�re^����������b��2t��� �i��M}�(sv�B6c_Y��:���7�?Y�xM�)�P�e%�2u���4�R�/�-�T�o���X�6���\7z����V�؁�h� K�A�&�(���^�a3ϵl+�����*��g r6=� �Љ�`��gk�ٞ��s�eG��#&�x���*��5õ��;|�����\��js}n��ix��������!��N�?������"�gw��yv��؀��L�Y].`�d�t����Wzan��>����^g�}q]^	�p�������4@�9S�<��B>���AM�T��]����G��u�間�":;%D�D�I{$m�HE$yJ��C,h/y�g:x�;p<�t���X�d�0��H��P��eRV^�Y��-�e�?%#����ȳI���Ч�A��o�t��lo��s�צ�t��f�7d�R�A��kXM�CJj�^]Jzk�HyR���K�0�(\�ob��T4�x���,n@���1#������a&{������e;�n��m�ە&DΞ\�/�~~Y�Q%���{Y�M����y���g l�wi%Y  !������@�tN����G��V�Y/e��"�hP�픍�9��u�ǂ��>�~�,�v�y<r��+:l,�J�7( k�J/���	�?�'xT��G�*l�+=A˕�
b���Q�H||��'���f�6?��,G#l�)����ziy�Q؃^�}�7��� ���-�ۿ�Z�������`�4G�Ol�� ������V2�#`����UN:fI�{F���6J,����>�h��.1C��w�*U��@z������8_�k��H�Z�bq,�xJ߼�9��,��A�}1LX֠Xsz����o�H��tX���6���&M�oY6@p��o�V�
g�06v��"B�g�s@��h��)us�};��-VO�
�l�h��]3�n�$|�}�G��E��[�X"SL�< J'���`�ӕڛʳ!��:V��Gs�։xz&�䍲���dPB��D�H|�0Zɽ�"|�X�x���˅�N��t�����c�t���G�7�$�g,�JW�X=�n���AvZsb���5�
�so���+�߮�.����z�@��~�Y*�����#�l@=0�]���� ��tpTM{�����5�,Z�V�m{+:�YK�?ݨ(_���;��w���#��M�������1�H�S<E���~�V:�w�!�G�C@�����K��c�4��8؅2�3�MѤ�xr/u+T�*��,W���5F{�H��Hn��7��TR��!�XZČ����I��n��@��=i������ژ�f��¨�3���~`=Y&���6(�
�������Q~���9��ֿ�%�x?b!9�f?n����`(٬x [5Ϡ2ە(H����`����Ya��$��Mن2o���?��  ƚ#�֫e��[m2�]}�}�#�(��Q͛'=�)�-�����#������!9���箯l�p���\`�쐵Z�)���A�� �U?�w(�!��ĳ(�����"uԬ8n"O�6��2��uг>��5�+IY~V��heE�A�,Ic�"q&A�rCM��<hU���{�c��:u��H9I��(SAU{�r��3�	6��������8��î]q��bZ��C_Yz�c���6�����>�a2�
��)L���I�-��_��4����Ež�+���B�E�I�+�;�~?�l�Xt�R�\�d��]���fc��:^���?��'n�Ќ~�V�ˀ ������1`�Z�@�ŒM�&�.�����dH0��W���e|f����<��.���t�<���b��F�K����R,�mb�G�I�=�rr����D'j�K[ߊ���n��9]��~<���l�1���>�W ��N@5j�w穂��oR,����~�%�w��kc�NF�.�=��j�j��3O}5b��cm�g��Qz�Ĩu�%!mv�p4r�ƣ��Nf?�Sn3K���x���Ci�����o4�ߠSa0�ݣYH,�_Q�~��mn?�2�G��+"�$�;�7�7۸��@�E��s��7T#R��&l�p4�t��=m@�&�����S���� ;��gl��4�dn�<5x	v�r\�*=|H�>5�T��]�ڟ=����ׯ`;qփ�$���?�	f�W/���z/<@�8�寉��G�O��ڱB5)���SIE��4��q]��U�W|��Ō=SG��
5�h*?eSOR�̥R�M�uS`]���Pw ׻�Հ����3�;���9V����Be^�M�"� ZT}�j�p6e���E2޲D�s�i���VZE�o����G�	x�4�Ԝ`g�+�P�P�,�o,�q��f��Y5�aF�i6�������y�LB��`��Viq��JT��!��pv�����R
�)h��&7J�����EQ�Éi5�s��+˞l	8'�n Yv��?͗f�����PN�\�oH%���ߪ,�(ś���!�������S�-i�0B�:;3��Q��Y��T��
ݾw��"w���v��~�SI�̦+�L���yY}\�����I_~�Wf�Wr�	��}qx�A���< k� ���X\��|h�Hg�ٍ�J���Q��7�*�mA�;�(�>�<�UL_cG���
�8��;��+F3\3Db ��D�Z'w<���}?�X6�I�Dsä�`;[ZF�>@_�Ø���]<���ʑ�JF��x����z3�������3�]�M��$&:>�et�A�k�}���`zJ�g�����j=<��`
�8����:��x�f�|#��@��+8���׏�FJ�l�V�lm���l�x�\��"�
�a�\�}5�]���cHD�2ψ(K�̌+�]�`��/�i2�^���&Y�a��c[�V��!�2�W6��mI�tR����J�M�!K�]������j}�ܫ��V�s�)��&3e�\���F�헔�G�O�7��`$kL��J��I`th�Md��#����q��9M�	\�5�9;?��O����Ʒ���<��[�"�"��B�|QVhN=H�b��2ˋx�f�������h�)"= ��u*���}�����i�̐703<g�#7���8Ѥ����}���bY�]!C�N��]W/\�T*�M�pf6��ņEF�O�7-�9��G�J���0�ԫ�W�o!|��Ie����α���G�l剋z�O�F��ｵ���QQ��c��E���2lh�Q�?�2�?���nmyz��t�"bRr�w�⥗���|"Z���>i~����e���)�����3c��g�m��0B������$�i�$�:�0E����˞:�y�1!4�\��z���� �?��X��
�j�1 #1Q��T �[@v�%�_�V!�ľwf=l����m �yL �<�w�4_�1!�*p�q�1��9d�.b�|�ȵ:�K��� ��>����$ ��cʰ�b��P#=m���?���u����T�Ջ "(��D��c��X�I1��3���`�O>���@��:]������\��}�T�"�@�<r|��oz���(,^��Og�a#r�1My'�s_���u�x�ʶ���(�)jخ�8����K���3�g:�\��3�k�Xh{���e��pN7�xG��ulJ7S�@ ��S���w��Y57ៀ�2���E��³�)<����.
B&ˋr@���̴�~��J3�@����x���>�ҡ>�]��v]-M �ş��1z3lxl�j�Ìĸ�y��IќjZ���n0��\�z���FN䉖��v=�B� �ϗ�`�u��Y>��lȧm�#R�`���ԄP�b��1�����e593��ݮ� o����{��J�c���������O�:��4���ey�SA^�"Г����:������Df�B,4���4*����
�c�uu�u� �~B,���Cˎ���r����/:_�mxv��(��*�,P�C��vB̘������'���]<M�I�qv�|��Ӣ��WD�:�9V�(�Ƌ�$SR�n7Y�d�i���!�0���8�5�g�H��^h�����4��7�u�(7��J�x�h��3)��}�'�>g&A�<m�%�8�A�U�C���Z$u?���PɧZ/�֔�;�:��*���WCkJI�����e:�V��]0��9�:�7�Y��4fa��هv淹"�#��Jp��27>'?8��hS����c�J�0}�41�P̷qnߩ�/��P�'G��C�?˲�����}P�k-��4HE&n�Uڞ�G���	:_x�,01�E�-l��:��j^�}��?������W�_�ؤ?'�:�c�+�E`�?{�����)��@��9�J��ii����{ʹ�*C�`�fi���AT{���3���~	�\�=Sl�,��8�\�Pc+oRJ��eT+_w���:\���h�=���L��?ΤNݴDM	��K�@�9�ZhN��lH?"���x��$�d�2����_���
?�ᄃH����G���<��p��5�C;��j`�=U���eD�����t�|���@��R������:�`��.H��Qm��7yWX:��.��D���*;�g5-o��Sl���H:`��ߔtg��!��� <J�l�K�d���1pi�*1eOf���"�zg�Pj���3�M�0�u������E}T�����/���&H���u���hi�'�,��	l>���ǐc��i��EV5�@j"D�o ^n	��{���NR�4�(m����d��'}<m����q*�D���瓙��s��b�7�1$؊j�S^����a	�/�v|����"Rj<�=�m�����Qx�Zi��@��íױ� `������Y��X��Ѧ�4JTYG	s��?Mn&��~�z��@|录K?QnO�S���ڽ[��gB|r�z/�A�:���������1�hhR�1\NrR��f����Rp+<�a��?ߣ��e>������
X��+N���l�>j��Ej����� �I�Wz�DOhˏ�r�?ȯ�<ޚ�Ȩ�L/��̂�g�G��V2���D�(2!p~��`m��/�X��^�n�GG�
��9;�Mo`J���&{
������ ��i�l��Xf�Wɜl����*myjY�Y#o#�m�·�����c�{������P&*��h��qH�1��V��`��\� �l�?���F��Z�:��&dү§��>;�?%M�3���*C�1d���<���+O�$<�����6�������!,�~I�)����f�����y�t���m>h��YOK�,�EjU%�~�y36Kβ�g-�C��-爐�ؚ¹����~����[B;%SJI����߽���*�E�O��p�=�R�Q���@I-}�{��u.�D0��#�D��[)�&µ-_�R���3�� ��7E˙I�L��,LcLP4 xo� \��߱2����`���s�HP�L>�,I��Ѯ��f�^��r��g�RH&��`W�	|��ڰ��.�h+����τ�e�[���Y@C�tdYP���u��h��i�dH��vN���}W��1���؉D���{"ko�M�������H=��
YP�	%��o�l�4�AW�s��ȣr���c��l�BY�&i�#!�p�0��9w���)i�]M���N��ֽN�AÂH������t�;LlO{+w�7I�s@,�M�
�Z~H���Tq?����c5M_85���DQ��7ө�w��RТ:j��h�����}���ѱ��f���&t���f\���-��A��ar1�!���U���:!�NSm���bj�Nӊ�.WdL3��Ǽ����>�. v�.�����g{-��U�Β�-'k���!�+�75	j�0dR(J$|�]�I� ��5QuV�+c�e����R���W1�x+S�O���1̣֢��e��L��N��;J"��mg�0(�\��0c�zZ�$T'�yH�O�졯3.��F���_9N^=	�Z��T�����\�r��$���}�I��;�K����M��5�<��|����W�� Rol,3�K�s��C�`�~�KSz���'�AǖRE�p��.Cxo�,& ���lzPN9Er�r���ϖ_��D^a�U�ad� ��XKqp���ō�x�ln��7>GPW��	]���8����$Nz�gh{�Hx>��u���n��pM\z�ĵ=*ľ�*��Vv�5:N��B�5z���V���r���f�ʹ���ǅ���8oaCԑ�иޮ&��ϴSG7T%O%�r�O@֚yӛ�X;߄3ҏ�-.���$s# �R���u�^��N���M3�>a\[�I��;����!��dS���2+��~?Mڔ��`(������w�i��߾Mv�'#/!�衲��^�w��S��q�@Hb+0Ai��w};��$78��|�Ʊ��*�N��D�Cm|	Ӕ`��@�8��J�R�z9�U�ND�aF���Wۡ����j��(lQG���u�/y��TT��r����k�v���w���!Bu��x0B�����c} ��7V��㓃ET����J�`��L�C�F�r1\���a1XGpd�g�(��J��L�+ ��,�%0�ɵLOZ�kBu�b���[{}@�����w\�Z!ĚJQ�����W��2�b@hR���w����-� �?�������{d�T�ل)P���UM�=��7dR)��}��A�\!����h�z�ƌC;�:hso.�,�
0�����.Pޓ�~�Cq����������<p���;���|���H�ţ��L"�*31&5�=&fpV�ٗ�v�&m���>~���#�	���v�~a�?�*ݰz�l�i$	�߿.�n�]%R��L%g���K�fE�sE@�\�Bh��ݔC��q��-iI��lw�ޥ�\����7lU����+�	 \�Խ|���e�E3��ךX���r�^�'Z��G{��ξ��$�	���`�N|bA?���NU�M�1~ZZ�p=�1P.�Yl�����0(wS��r�!?FzR>Z%3dA�!$x�	!a�j<
�k���#��Xc63����n�wJ޿�͙����~��s����F�3~	V�&�n�J��ﭛ돕�O���碌��X���E;QUC�;#F΄��}[v�N���E6���9� ����]E��Ts0��(��̖V[3��b"i��\��+���8�TbBc$_qǼ�)!#�0u�0w�Ba���첌c��O��0tT��i(�����h�ِ.�R�)yi%+L��/�/���S�.�p��S��(E�q�ʱ�F��ޙ�+�d�S#��-�%q��i9�E�	���"��KQ��*���+�$�*ջ���,qL��j���4M�pLh�Z��~-D��k� ��O�����\$����I��"�Ԍ�%�!%-�⎲�w=�a�M��������+��d�alhv�oz�T���!�1�ذU�����}��b�����,�B�:a$//$Bs���s �I9�^�< ��})��\"����K�š>UTi���׼�L�)/L&�M�f_�.�ʫ��V.�q�(d�v�q�|���i��@� ��d{(�����Wm$���^	_hU��0s3$d�ZF7���Ö����!�_O1袣 )A#J�6��U1�ǿs�RkT�&�(�t4�0�5��iq�D��p(�ǯ�K �ܛ��Z�=��$���d<a�=[��tKC�����B����l��󢘳�T�b���g@[�?��hk�V�n)��	#p�uJ���Y�l�ł�k^�B�[����Lz��1�O\��)k�q(��ֻ���G��݇M��If.��sp=O-MV������F@�M�n:?��&�t����QA(S6��2�Ԩ�|Cc s����uT%د=�Y��Z]7=+�t���4�\�d�擘l �+-rwj��(� ������@ɕ*��2�d��!��mR�ex(� D�.2-d�;�3�c��
�G��FR I�1�D����쀅��)�̘������?���|D���N ?��d�8�:��Ͳ�r�h2Q��W�ö麝£[������6��UVV- �0�T�S�9j9�`V��S'qΒ�N���P� 31��qq�1�� ��b�Bs'�\½)���pxH��p�j�9{�H�pE	\P}"3��&�$���@Km%aSd�1�V��t��mW�����;uJ�(b�����#��& ��x����OH�Uɯ2�!���17�ra�O�����Fv�Л�F�.��q���
�ª����5?@w8j��?�D��tv}�j�Y^8E�J��	RZ��Z/T���O�)D��b �HB9Z'�͘�G	���Ëi����^-�4��
��ӽ׭<+V�^�K�d�p�=d�*Q�(��^�w8����WF��8�H�/p4=ęzm���,���]�"�\�D�2u�C1G�L�n ����5�s�|3��0b�G����dg�B�~����KJUKX���	�	`	��jc�>J����,T�t�|@J�3�+.�L1�PB���☈���Lvx�:q��8�UB�Z���1bѡ�ޡ��
�g��!������3�<8�{�:�Y�����+o�ư����$vu� ����Az���5}��T?�[Z:��5��lJ��Z��:�F��V�2�ˉ-��W�'�ϲĄ����Ф�Q��\+�m��P[��6�^)UψKI�4���b���,��W����9��҈��� �q�O�������GY;�P��Y�_f�p���L?�/A^�ƶW{�i���o��&� ���&Cd+iZ��"i.>g�f<�w���K���㭷;�cĦ&q�
���@���(t�H.yN��p��ne,V/fs� �v�(j�4�B�VJX;vy�\~_|�u��,T1X6@M�������"�9����q-1�^�w�����7"���K���-�,�WfE��uu��J$���_p";�V�[;�G���,v�׻D�x��a~���ا��j�I3���jy������������B�@d������ܵ�+�20�/��i"�'�&�<BD���s�j����笋>l�����\����`ע�b�u��)�8a%t��7�}-�h3�M[
���� ����<{�������$�3��o��7�N�>Üi���>f�BElǚO�Rhbf�%9��DC=�7j�^���%�`�"ɁN
�-��Ѿ��(�����[���"�RN��b�\��D:FM���:�n�6���L�8%f[!�wO9�|n3ŵJ��j���f���� �Q�Hٔ�$EjQ[��R�d�i4�����eL�=3��V�?�����G�yY�Yg�c��|Lo	Fx߰�����//L�E���0u"�:�J��üɦ��'(����]�uRjv�wtb�>���t��~�gy1.���_���'±��v�bg���RK���23O��[3���W7�}"�*�I�
b}?)�X�;�a�٫�U�"��5����-�:S
7��6��Ц\���3�8Q[���D�l[� �; �.�򃢒�%�ʃ^�����Qx
QCߟI)���V<o�l���#dB�?�Q������:��2�P/�>�ݮ�R�q:/��&?Đ��u�T���vZ�H[32O�+ʸ�;@k�G$�0>j��@\ngx�ef�#Z6��v���Y�����T�x�Z>�O�8ǙH�/d��w(��u�&�#�
ǉs�|�필1i����g)��r~ ���{O��R�������j�r$����_�G7ٺ
+���M�)ܠ��s;x]�]��]8�حvo���8_=�0���-�[� ����N5[Y�;(nq�ؑ�l���	�Hp'&�������H�Bʈ�zF�FȊ��t�z-��Z���h�&�	+��L��"RTv\}u 4o��0����>v����L� �dC��;�x�^�߼x&%����J^��6���i���%g9_��sGې�/-��
T<E���\c����CQ��r"���(T�,+Ҭ.�����kB4��!yW([�]�Uf%�������c3O��hh{1�l��"r��K���q)�g��Na���[��ĝr�W��qS�d�
��RR!�F��^nv4��Y��δOQHT��⍺�n��J�&��,�nQ�hC�\L��`㧒f�on����=2f$���u�C@��W��@se"a<>�^�q�_H���i�'�zVF����lK0x ���� (E�]�dKq�`b�I���_����������/a۸�?E�O�URV=���Zp�be.���#�H��>%�#¥�(H,`6|.u��RP���ˡF�?=�w��H�[����8B�Ywy0K�p���׋mr������b�g}�lf�4�δ���s/d[#[�.��������-�+�ϳ7���Q[g�lT��>7%���w1H2�?lƂX�G��1���M��� �|���w˭�����E�Q�'��w�7���mϟ9L$@��dk�yU�`�Cr`�y��o�
���u��0�O֩�����!`�T��ig��$@lj��BM���%l�Y�@��4j�*���g�}v�&�4"Y�o	`ǅ,��t���c���|t���An�iJ
��2V����*��&�V����F=�A4����@��+Y�V����h����<�}�T��z�<؛j��'c`�<�l�sr�|��gW�w�|�d
���U�� Y�9�i�l�R�� k4Uv#['<����9��/�,�������K�Ob�_�}UC�{�I�e�*
�L�a�t
&��rOb��"}6����״fדY�䚹zv��C�O�T�[J^<�v��foeSV�lw��*�7+�X�hL�c~�oyfE!4�8Zq���-�N��)#��S��v�(�ٌ�V�����*-R,!�|}˦��[����Aζ�u���J�_\k��^�q��EO����84����vN�@�LC��M#��ƣ���xe]:$d2|�*a�Oݝ��������a��ãbYE%Z��a�p�5�$��=5��,A��']�	��J�M��G�61?��T(��"�u5�q5)Q=�.`r?V��+���&mhݐ)���I�&��	t��K���0z�;�uއ*�(�&_�d�f��홧`��Cg�;3�
�M;'�A�l����U�6�=�@�$�뺉���qEv*�[�6�Kw�'��,��Y��
Xc='P(��S9��.��[L��i��EN��m��I��9��;�%��B�F0}����Y�����[mK�q�����+;*��W%_�T��6��<������[$���W�*��}'�"ۃ4ۺ w�J�.׳��&��w�WLëOz���$��,�v4���g�Y<

��+8 ��̚0�Y+%����nL�	"��+������p�ߺczQLM�nfޟ���S�z�
�fO��0����i{Eڍ�ӓQ�^��-�$]�(���5�����l�10��=B��JA��v��.�-���,K�5�<rW(�K����h��;���ʍ��z3�`����s1Y��TQHIi)\�F8Yl���M^gC��[m��=��%8<���z�@���z��D�˽x�<NOy��$�k�j���7�
���T���JK��^�n���	� ��B-h��΋�6b��/k�O~��o�nC�K����1�_�m��"wfٿf�mz, �n�B䫼�g3�����V0 ~��-og�z;�y�^���%ܿB�HZ��F�(+jŠo۔�5��Z���>�xd
#��8�t��{Pw8��|��>V���z�=7��,�t����Y�t�,Јk�������E2��nP�P܌J�4F.���߷����������~$����_�Xr-��Q�9e:=�ؠ<G2(6\���o����)��a;��(�Nz���z ���e ��:�!=ݠR�lm��Q�l*�U���o��w�I�*L��!}��m�C4�5�r�A�9:��Z���wGg�e��=IOB�d��6j�1�����`���|���`ͤ�!QLܣ �G44\���&���s���e@�]�^�/>Xg��a ��a���?�6&L�s����2&��~���Li��=�l9�1���) �3j�G���� �Y�>D�t��z�U)Z�ń�?�o6�K�{��� ����L��a>� ���:d���$(T�����5 k���CfG� [N(y���z%c.[���H�wk�`f�F����(�{=�4H�;֎i��I�P�>��y�e*��ؑ�O����h.�O�K˶yQ��z7|?��ą͟'�x�Xo˖q �$�;V�.ZItQ�\���=	��_<"T�*�ϧ1�Z����<,ol��j�~km�qi:�J��8�E��&@�����c_%�J�:���PY��AM��`�m�.��6��Per(�*�I-���ր(,�]?�%}���Y#�:���\��پ��^�|yD�6؜����HHV��eϑ$zj*���C���"��N�6؟�/`��B(��#:\�ݼ.�J���U�te4)������8� N�5>7�(�D��.߈��"�בm0��* 6B;��ǩ�2C�ŷ�i������Qe�Q܆��[���g�<��>+�9���r�3��no�kMgb��M<���PP�٩e���迩=���d����C]�g:Y��r2�t��w(o��NW�VH}��*}��e}�����}��͹��Q�
+c�F���6g���)�/�1I��Y�-�`����,�W�e̠sd51m���Wjr�=�l�<��|ݯsM��(7��k,,
�J�M"���F�d�_�N�����-w(T�j	�j��4�ʑ�4��������_��{�Cn�4��4R�8�^$��?�5������a��䛠�����b;�Pp��̔ .lo}�7��W�(I>rz^>Z�����i��a8?$3��Hv/O-S�T�̊ӈs�wF���fN߰ОX�R)���{ p��!�x�`A��5�]������0�i�,������jm����v���U�i5�lh[=bѱxG��D!*.y�W~����Cde��%D��2,ny|��8�Ϳ����8�0�^Z��Z�}��_OŅ��-�W���_p����j���
<9͕����h;ZQ 7Y�,׳Dbf-��!�W����
	��P0�L�@8rƽBl�/�bߖ���+�V;���C��b��0�ζ�rA��B��X|CV9��y�C
n��=�.��'I�S�9#��Q)�
���������$:�.��M���T�'s�����v}Sܔ��Db=��� ㈥�D��,HeC`��jr�xIw��_���������/d��)�$&P����E/.��_ЗA[a�U�����ͭ��v<�/k�f�9��#���1U��a=�@��?Bm~ߒW��h>�+O0�-(���T���k��y��@�����,\)�X�31�^5����57���b	K�m�˟�15���~��ZQ��SϤ�|7X���P����`>.�$i�����x�z"\nW|��$�7g����Î�=Գ�� e�����, �� �j8y'|{���Drz��9+GB��ĦX��ёƩ$�^�y.�ɒi�y�["��o9vW��ž������m)-���Z��Bo�yےC`k�i���h�Fiu�����-�2����x�˶�Դ��}+���奥�>�:N��Ǻ�dz�W[���F�Y�%,=I� �̚&T��@F�B�(��x����\%�"� ��Sna�vx�:����|��:�#��ý���E�#z׼*���8�M� ���)5KS|��ןPW����@��>�0q�S��f+"�ԑ����1+�r�N��}#h
����c{��ډ݋l]�X����<N�;�A�/�@��)�9���ՖU�:k��;��l�6��n���K��Ȟ*�7~$6�����籫��G��j=�'��Q�薷��I��Њ�N)���W��!!���\=U�m�>��8Zԗ@�y���-i\�
I�ln�� �[�G�-͘$�c��]0p�*=��z
䐆ζ`�Pm��a�2M?B�SP]�Cg!þ�D_�H1��ោ3π�ûR���3��MW<�D��z�����R|�5����g���0)���N:���S]F������~�ڵ4�0�> ����nˬ����<R���Z0Io�B%����������G�4�|k�V�B�&-g!�|��ԇt��X���fs��l�a����WNl�X��-^�'?�!<�ȿ���^Y�Q�k5����L�Yo5I�%���/0�1��/n��p]b��(IM^���$��OҼ+��O8�0n��i�?������:2�� �8�k��y5
�gu�/�4���=��-t�����!����e��ݵ�b�;K��ğ�g]AӬ�� �}0�h��ф� ��e�Ay{f5�"�`ع�ہlM���Ƹ�"�-J��qH0��2@f:^+c৻�0��K"/�� H��1�y'S_��A_�r�|�2U��gO��t�|$��8s\������'�i�s�Gc@���t�~2�9�Ra�j�~E١>�i�����j]�9N�/:�����*�X�<\_F�V3s�wE��Ge6X.�j��^󿏙pƇ׫�`8������tC}k샪qiN�jtPI�W��T�4!a��y��ѩ\�a4�v\k����mc�!�X];]���q�bYā�4��R��˃��,n'�K��nT��.�\8My�m���X�J�<P�{9&��(�R��z��Y.�~nf �Q����ryy�U� Z._i�%Q/Ϳ��lg]�l�XϷ��Zj̮@�]\e��%����_�AA��r!u�;��Tᮙ�(�Ѷc�/��:"L_�&˂vB@�߽��,-�W��������5��vG/Moj��E�_�~GP:z�
j�CjJ��<�����iG��%�]���ͷ�O��cx�M��v�I�Ԣ�.�UTN�f8���@ؚ@olr�oR�2���]]�����g��f�X����),�v���)<��	��5����R{�oq�{��6���im#e�Q�>�SW�� ~���M�����̯[.#}C2G�B2�WF�[�L��A]�]b��q��9\GJ���|�p��&v�ّt��ޟc^%�[��aS�Q�Һ�_�|q� �tAM-Kֶk���}�[��#���(������˚��XH@��l\��	@���.�ay>�+�B�����؟�B��wk0��@�w �"=�ZxN���ނ�y3�q��F�*L�R��5�㛐 ݎ(��Z�H|�`EJt�"_Z�̶ۭ7F����8���{wR�L��3����#A�={�c�p��JM^�A)u6�p���Ӿ�� Z�p]5A��zv��lG��ĔQ�5o��T5�'�5��5E#�QuFI�"�K���rPn=*>��
�#-\`V��ZP�����	_�1|ǘ�H�;��Oᛗ��dX "���E��D���P��,Ю��r�W
�(��X�Gr�6��4�.��妽��X�M��Lrg�ڼ�)�I��Ʊ��>}��Rw��X<�y�^��i�������
�;��AS=��tK]5Z$���a��%@(�4Rr�J��A�%Y��d7��9M�':ts�d�v�l)9.�d,��O�*���CbKY+^7��m�&^�Th9���W�o@툖\X�}�8
r��ۇ{��3uA}@��Vfl���C.�������Y��{$�O�� �Jk��$r����zl��V�{�Q��AEt'�����q�կ�S�UεM\G��m�\���BMs:0�Q�^����!Ze���H��P���/��p]��4B[�ױ� �*�-e���{He��8��[��Si=�eQ{�[>��B&o�ߣ�G��$��M E�X�Qf�Fܘ�0J��{�@�P���}��d݄=��m��ȿ������H�Gt+�EH�/�|�['(e���Q>���th�=-V�#��}�DC-��_��kۗ�ž�*�X0V�P�,!�Й"u�ߤKU �����j��rＩ���m��꟫�M[��9�����e�lZ�sG�^W����~(���?]1��Ȏ�8������9�!&"�%����~�H(d���j� 2�J�O��B$�#y�pn��Kp*���bG�z�h;�ӿ����J���L�<���肕܄��.^Z����MU�����bY�L�EphK���>�iȣ[�h��z��F&K��-|*�Ώ�'��T�±/)I��o�}:��d��R|�٦b-l�<���l��Z�`����u��-k`�z���2/�K
��?���}WA���>B�#�,M��8j�W��or3�p~^b�F��dm��C����Z�F��������V`��\ܥ����_>Dc�zoA��P� �����wn}�V<�� �P��t�^��.��l��`�.^&�p�,S��Q����ȯ�ϩ�O�s�L���f��>�s�Ef�K�p���`����m杰	��7�����SITxi�׋Q�>/Ǳ�!V���6�7���9d۪H0�4�lj*ڬu��'p���k��[�Vo�'
�Ҿ#�t_��7�"��a�-��|9����oz,��K����e���e�|I�:�⋼8���)��Ĩq#�8��qkS/��0	S<OZ�k��O=z�
,.�pQ�e����X,(�5����Y��tE�#��dެ���>���՚�y��咠?�oX��P<*��f��G�¹�U������Y۹A�$��x1`DP��=��c$ y���Ĕd
��x��gǺ�" �9E�0q�	�X]��J�ɀ�fdJ ��+"UI	�C��=Zku
8���&;x���9���pЃxن�z
�A����Y�|�Z3�J"��<%��� ?��4�P�5	���)*M��o���{Uzn���1SiB��A��oL>3����I�h������,�bM������>^�%�h�������<�Y �U�W�&�v�ͩ�g}��'��N��e㗩GNe���$}�4_��9䴯(�œM��}�i�Z鎡SwuI�~o��.�J�����י���2��bq��b�G0Ы-p۝�ɦSL��yո=S�
o\���:���8X_��U�6�as�fݭ���4���2㴆Y2ty���X�~0��t{��Lq[2�耙����ӷ���o{:��h3������MWags��9��5����=n}�U��dm�� �Ʈ��b1�!<��@B�q���:���x�xMm~�?U9����7�7H�p��9��H��g#٩�;�����{#��^�c�k1fD��週O��5�����E���#��� %���B�
ٯ�]��B+�r����|����6A��c:�,��0��o�cx���qD �|�g���ta��STd!��(<+j 'G\'O`���O�?��)�S�6;q	�*��fY����R���s�Cɓİ��N�Y�w'�gn1$�,��K��, �19�zKh���Ș?='��HN ����df��S.��P~�t$څ]�NU�j��k7B���A��Em��41��Ӹ9�%��I�:��t-�H��lV���+֓�S	O�GOW�����#�!��M�~@WVGC��x�v����-������*��$��w!b���R�r�d�K��d!$b��f[�}C��7�ӱ��W�}L]$�/�@V�u��؍¿B�[���F��w�ws��G�2���h� ���*Z ���<Y3?����|kW�R񨆆O'��!��s��ɒ0-HT��l�*�.�}b�(�i\�_W�;�kh �O�Ԭ��c�W^JrZw9��j&�G���?���S1d��|�YY ��8[��V�dYtb��VD��0���#�a��-������R����OJ�H#E�TH�e�r���'����"��Cݍ!`B��=���bA�z�u�
$������3�������9���J��НG�On�$\�0�@�A���#�~��y�j��8]b+ ��������
Jҿ;տOA�x0�bNl�X��(	��E��n�[e�C��VgS"�L\��*�sO]�#�<����ԍF9k�Luͤ��6������=��a��Ϻg,B*U�]���0��)i셺�6�3��lO�_��L��
���3�,ms��Zl��YX�D��Y��:����F�|�?0�wJҥ���cBS.#��m���;���^�7鏍2!�ɢ�W�Q��N����8����G������e(�v�=I��6-�Ce��dn��<�|C�=To��e�,#�N�p���qʊ������,+��)m��&���D[w�^MF����V��Et&"�������:�����R�����c����av��Q��:��}V5�����\�E��/w{��P�ny�5�������
CX)M��-�S����������V�Юp���N� �0�W���fL,�a�)��/X0jp������b����dP����*/r����Ѡ�g,����Rr�s�Y�S���l|�������)ե��jjs�q�3����I��){�Ӯ�1�q��m��^�W�A��mi��sl��R1����ܬa�76��ì.5�c���F�Н��=�8�����9aH������0��},���G*B��2��P�(�¾���ؔ��JpEo��RSK*<�0��%��.q	=�<j��~�f��(���*{�#��8���to��+��[���}�َ��-F�4�.�]��N�U�;�kY���R x�:bI-�!g$��눨����%�߮�� ꕌ�V�N�x��Y����*��PE� ��)�f�763JY,��JÉSPEY��Evnui�3�%�2�FZ��	�h0�y����%?�;���)ߣv,!�	�s����_�*�U`�䦎�9�+�B���H��Y_Wꦝ��[3IGR���k��kQIQ��<�~B^H��h�
�1������.�S�I6�N85��myQ��v.N�I�Ys���yB�u	�ھ��~]lio��MJ�(���ǒ���Ab!��٠����S���GE�� 4�����<eYya?:=x0�YMH�#�È0��Әbĥ �Y�,�n��9�ш��%:a���ܳ;H%�V����*H�M���JÐXP���hş���^�
(b\Tb0��(<�=��fݔ[#p+=�u��F�gN�Q��� Kk��oB�][	%x^�k��WX_�݃E�!�!w�(���l/�&;��6k�W&��8���0n����:�0�l��e�Ux�{��ą v�d|Y��
8�w���?�-��m�Y��z�,~bZ�Gx$�y2�rmQ�ט�L`�)�i�����d~����z��DQ�G{�΍Af>�U��g;r���{u�ZњA��9�� ��HY�t�Rw��]��E�������E'/f���|[&�29��_��*ް�5�&���gw�Ɩ�++�6�;���P��Y�@D,[�JC����y̹��x���i_������eu���L�Z.���)1ӭ�:�7q!�1�(F�M���t��ڼ����)���f7;�_���g8��]�$��f�&��nԬ�N����9呪�)�`��&���J��r��|��*˻�+�ꄶ���}�Y�|�<����5�o�(Y{(Y	O�ߠ��[�[�_-t�8\,����b>�!���Q����/�R��S����:E�R2<����RK4}�APϋa�~��N�"��R�.x�uUR�d��F�ͣ��Lb�	�N2��>�L�f ���p�M�q�'l�G���b�Xǈ?�A�IQڇUd�$�ש7�P.���;���]��	h�RhX�����r��z<� OGө���h6v�P<�qT����ݠ���-�#��>�����Q���lQ�)�X0wOs��Ұ֥�_��o��\e�ܟkD�|���Cl����>�:^2TD���q�o�
�b%[)��4yGòzw�W��|]��m��
���*l;6z��l:�^�.yنWk~5�v��M�=T/�/�u���-|�9��8�Rsq:b���a�|�kQ�R?/�?	x�H�k��y#>��7�#F�s��*�~⺦v�sW#�w���ˌpߖ�5���:��2�g��T�Q�=v��6(�@_���H��0�Ι�th`����ۿ
�[��K��v�i��6w+�J���m��3K��$c�
KO%��+�N~@��:)���*y�p�A0|~�E��K��J��c����q����d�^P?��u����e�oY�YD�/�(�ϲ�("n���?5]5M;;<�/'�RثR,�&"�!�|�8�s��p/^*���TK;�w����-�*_|� ������^b[�Q��Ư����k.߲jq�k��7�Ƽ�sT�Z%1���]F��G�Kt�6�
ڥ�ţ�������e���܆ӭD���҆;+�����-��V��3��@�O9	��3������r;h�\ħS2����KIl�ĝ���}�NRyOė"���y媴\�S�/�˷@�Ϙi�Tʺ�\�W3f��N ��Wjr���@a��Ү5���s�% ��	gq�<1���&��/Qy3
�b6�!n2��5d���iu��0Լs;`�؃t	"�l���������gcNj�!���Pׅt�E�Xz����ʍ�Eǂ�K��z�e�J�3r�#��'�ƺ���n�hC�3��B(�Mc2lX]�1=�W����H�v�Ρ��ӳ�԰"^k�۽�K�����;�	�7��2�{O��!p?�����n{,ʥ����p����_�a�N5I��k�cK0�[EM�=��I;�x��Ii�}�����+�c�x^�Wy�<x��O%����UL�_bd��%�«ҧ�Yae�:��&�Y,������|a<�0FY�J��R���]���Wž7-4��l6�U�O`�a��a#�N�v<Ն@�4H.��[`�#C�b��c';�gy�/K�V���)E�NE�����h����6vU"t�bSQ�Y��ĵ�f0-r�~�j��ɞ2)�~�	���sz�>�O�+*�2���}fu��>�_(�1�����(<���N��ߊ������|�%ً�k��o��r�͊�h�uxޱ��?��jw���X�3���p�L�o�8��W�� �^;ۙ��kk�'�B�#��>X�ٯڬ�a�*����|i�ō�פ�s���w��;+p�Nޟ� �E�1)#��������o{���W�Ы�=�ﭬ� ������d�nX��-�]
�����%a��#�=^%�⮳񠒤��]�����#��ٍvC�۷��*�;n�����`�Z8�0lF����
�ES��8�)^B�����8�����Sȑ��0�s��������В��Y1�� ��q��^<��v�Z���0n����f��܂�(mn\�։*J��Ś¼��|1BL&J�0N&��k	���/�i�m���!h�;(p���AVzܔ��jZel}�C*B�i4�*yŗ�t$m��,P��>VIѓ������OK����e �U5FQ�f�D�w�%�e��eN׬��`�\,}�`i�����U��x|��Z�!�n*K��9��!�&}�����d϶�ln%U")Z���ЃB�iWC]��i����r���jŚ��) J��,��
���/�G���DZ\w���80���*�k�[Kr3��*%]Js~����n�H��P�13�ȋ]�����ӷ	�x%��&�~I"�Ϡ��c\�Y]Tֱ��P{�g����������;�C����iaA~��s\�d�~Ju n��6D���0r���Ae���yu[���X���O��͇ܮy�VG�+�S��=��������q�ѻ�7K��,��p�|S���$��%�[�&�diE/P�8C�kȼ�{q`���w�j���$:G͙),��Qy���Ø��\ ������2��g>�{tB-����CO�!��KZYb���P�h��s�a�8GZW5��*�(�<5$��Ϟ�ֵ%�����[5��*�ܘ
��ͳ-IA����5�<��/��A�r� �ț�5� ��+�Z���3~櫨�Yy;m_$5���S�c�h%��(��i�{�AK��
���:��z��ܟ��S�U�z�{�!
���b��o��X�(��}��R�щ����H��]Uѿډz#�a@~���z#S�Ź^&�e�Gl������h m�u\�[���Qb���"���(gW#��S`��2�m�a&����=�ڜ��I� ��#�<3����U:�oZ�2�vvc��4��uaR�l \3�j��"��Zw��tc
�`)h�t�d�4�j�H�D�0��ߒߥK����r	5n��beX�������MY������,��NO��s�-InT����ވ�V��� ~fd�y�KZ�sV��GG0�|1��p�W~�[G������g3@V�d�Y�CG�����k��݊��s�l{��:�09��}k�Z���Z��C����H��&/�����>���ﶱu�<����z�c�2@�Z�=I�Q��n|��T�����<�k��J~(v\&���mN�/K��+F#�}��|ɯ��\Li5<b��� ���c�ݖL��p�{L��"�m*���	���0��5(���Pz��^=	Rdϝ8�c)����:)d���uP�܃x}�=��W#3Jt�7!�q=6J��zqv+��{�p����9����������`���Ԕ�m�>�,�E	����pv�{�oV ��d�(� �k�D�(i����_�͡�ñ�Fj�.Wi�S/���3�63Ls3[�Q�ꙕ��u ���(��لgJP��?���5e��o,JL:�i����Y:8!�N$4֨fe����%���ׁ�0^��,�VW��+f��)���K���q�-�A�e��O�4�MK����.��>e�K����hb��F��Ģ�%�4��3z�D�L,Ħ��@��?Z,W����M�<Mq��xf�@��X�S�Y�؂/l٨ZS��b��=A;��U�(ct��e�55�s��^��ެ����t�2%���Ǩ�xaՎ���8D�ס[����h�<��9�����Y��\,1S�_g21X.!ɸg�4��l�n�M�H`�uۧӼ��#�����0����"���{�>�a�o�N�w!.d�hO�b���*�H�TP8��`����?C����1g�q�$d����{���	w5���!BF��f��B �����-w�1��O-���P�B�c	�Z
�cǯ:�K�V��!�Ί�a2-����Dk���7��!�� i? �����^è�W�a 6��X}Y~�ng��S����εƢ)��[fVL^)	tߒ��y�c�>8��
`���p���#դ3R��Ԭ%�ԏ]W�4s�����V9Zm�~� 1!�ۨ+��o�;��xɱ����$jƳ-��y*-��>E+֜�����ŧWM��T�\s�/�F��bs�f�����\n8�[M�BX���q��b��+F���S�-.s3�+D�oZ�������%�S��r"�#���ИD�-�<N���9�z���<��P�>�k�����3T$�m�1�[�* ��v4z�0�#�X�<�e��3c�bX�D̥�鮒&h�BO�])���O�8�����L�:�z��|:�N��FD^ /�R�O9`��T5n�u�Z��_�l�=�P%cR�?Uep�uX�1�������)�Q4]���.��"%r�(gJ��碷�gy;���Wz:�!�T�
W}K�؃�c��TB=9p���ҁ�T>�mvZ�ξL�v�!�&��ZU��K��AC��!��J�p�U��˜�DZ=�q�Y�����m���P��U�����\"%Ɏ�M&��ʿ,�l����f3��\v������T��)d9�{�a�K��}<y5Y�ko˹�, K��(S���%I���!,�k���&�G�dҚ{�8��P��z}\�Q$Ҵ[�m�cU&��]3i)If�38]��7E��ր��A�"T��v�p��e��}�_)A����L�m�=g��_CǸ��vCV�}L�p��_��7�,���|��tT�ݙ����_뢔�M��#�������'�rq�[) hCMϦI�&��(�rb���h��8 a3{�f����)��eA[W��>�o����k�-$w�� �Εqd0�=��i썺>�P�� ��#���v^҄�2b�}j����<�7�
���r�~�-��I�ET߇�Dr��m%d}����a�����[m�U��]��H��zS�f�W�r���`e�Y�L�k۵� A1ׄ�C/�!�0��HWX���i??�QNؾ^&��/�9�6p�l�կ4��(���G����&�j`w}���<z��5��q�7qL� �b9�Ι��ŉ�:��0�G̷`��,?�F����ʡ��gB�`z��1�1��r:9��Bq�T5B�LҲA*�[�kj�A� �\6��\i�K�t[�+�(���1u�Xz��$��FS2%I9��5��U�����|�I��A}c�%C�L[����U��&/\�����@rd�%<OP��Lt|�����~/	���B��8'%�(i��n3WY1�ՓU���ߞ�6�_��d�z�z�&��v )#�ʃ�yB���}�_�|3���^h�7f���&kϙ��f��$�ߑMi1�z�}}�`oü��*��u���EG��rW��S�P0]eJ7���xۤC����-�<��׃���"�7˘�������ZA,�7Q�w��AB_\�I��������SEv��S��^����S�.�^�"�ԏ5�e�(���ƺ�yϱ̱۹�-�-��}Nx���?e~�f}K�Wx�9,��E�}��_:bG���q��8 ߰<'����c$��������0�����e�@���t�?�ĄTf��Z���9�NgfI>i؉u��/}p<i���ҭ�)\k^���� ��|��/����fIjx����a�Yit�nh7��7
����¸"AY��'�9�l]n�������A��ǥX��ɷ?sc
�6$.�����ѥ� �_�IEg:��_.˧��2�:��h���EF�r#���5'gQ�r����G��!���-����V�'�=<zƾx������z6�`�c<���F�����3���l1iG?��Y�J�4f!+(}/C��ipW1��iVpp.�+����8�C?�C\ma價�� �Pn�����d�d���7�O�\��v娇22��@]�>�q"�Ū�#l)�R��Q��������#�`��?���㗶�R%��gP�NI~�RB��U��bf�7`�o��:BJ��O���u��a�i=�4@w�P���z�$�ê{8+���Ptѵ��|jGT!7�'p��	L���u��.�*�9v��R�L!؎S�������M���3}�oVk���X�'<>��:���֛[Q�����B����W�H���d�Ԓ�U�V�����*����"i?�p:1cF�:��ı�k]G&��� j�VM{1{�$��_δZ�Ե=��ExO���Rg`=� *��������fe/&`�^҉�JUa�A&��� ۲���&�!����T Ƽ�ON�H~�+MA�*
���y�KG��<�Cy^{e� �_�"��P�ؕ��F�C�V�:}_���%��L{tz��!�ch07ZL݂�?�*i4�}GŦX��r�@+�w�.}��3 09��~�c$ ����*�������K��d�1gzi��Xc�������lU�L�����V&��^X6��Ĺ�
�VFF�;k��'	�@�t��P��v���Þ�&��"����?��D����w่<W��"�$���*� �� #����r��l��ɿuT|�E_MR-Y���������D����NU\f�0�g�g��dWT	q繽A�ր��of*������/W�L"���9 �j�F��Ǳ�g~zrx)r�$
�����j�b���ս	?�w�P�y�D	<�����0�f$٤�#p`N����t�?�)��[M�R �Y3T����}�6!�{b�$��/��Q�Ӎ���GB��",֓�k�?�Q���s��&��t�٢r� ͋h�������Ƀ�^~�Ō��۸�p߮�C5q��WVk��jyZ��geS�-�}��\�� ��ޑ�tC�Ʋ�09��g��m��4}���)8ʓd��K��;y�aZbr�0 ��EB�}ӽ�=�l�7p,-z�#�T��������+�gk�O��V�m�	~��ϥ���]�&��{\����#�&�����	�\�'�I������v�~�f�,��qM�5{�-�c����*� ��Uߖ�LقoVy[N������dY�ߑb1��mJ0A���2x$?��̂�zR���yk�`� YY'g�����x������֣��.+����=��5��uOS�t��gU/�a2�y1Q�kTM0Z��t�u8Z����6�;E�8�5T��"��
��f`�X(��ؠ�Aw�j�UǱ���6�����f���4�NX��iִQ9�SA^Aѩ|��`���a

�L���%��7�C^�Y]�n���{~}q���=�o�Gd���>�;�7,M�q�I^��j*���qڒ2v���N���3_R5L�8�Ѽh?[pO[	�+;�5���E��y֟(�i돽z����I�1akSw��R�6K|-�p���U��}�~����*�ۧ&���9���e�ru�����iq�-DD�:��D��C��r>} ���PWp߂�h�]�ȼ\�������A@}!�:́3���(گ�Οn]�-t��a,�c���{�p��(4kn�?l�X#���Ƞ�P���#�Jǲ�N��� ��9@BkC��nr�\<�P'FtbMU��ԱF�i���"[b�����0�b�A4�;�u��Q*ڴy��_@4�G�N2~?F�Q���p���(�|���@��>�N�v������>�B��u�B?3;C;Q3>�ڻ��}���J��k�m�q�����j�9��f���J�Ҍl�����
���:TU{~:�N�*?�Ы����G\o0��3 g9X�zg0�D>�C��^��㐨S[���s�6!8��2����D���(��{���x���E���yZp�	�<8�}�HS�g#	�7ls�^Q%��*�I}q��t�"Z_�4�	��W4�K�5Xr�(�=��~��k}�\l=�X�������!���;��>r��tzP�?l��������c�Z�Awj����z�(�Jƒ%E���21������d��8<�'�n�.��j�>�Wq��֣�O1ǩJ~�HH�� �����ݨ�7$��Q�5iCm����U�dp3Fh|AYGj.�d�c�W�Qn��A�3�@f�W�o�9\�wH���W_��q� ��@��3 �v~��ި�f�Vl���Y���%}�lN�3ÚQ��@rƭ���������Q�� k��E�����:���p�2����R��.�cÏ����T�X�F@a���I~C�c;����q5�pB;�C�cY������B��s躱��v�����I,X��3��s���(1׻�#��0�9���y��E�];��Z�B��r�l��c`X}M�.0����?�>����W]��MZbتO��'�ͨly&�,�àS݈������#OX�u V�G;�x��͝�T��E<+Nvٮ,�P��X���Y��иjө)9���T{R͎�u� ͋�}��=6�3�.p��ְ�{pz��������h�O%z�,��9��n�����B�� �[P :e��+��	��\Y�0~���&�-Zݱ�p_�� 7!ʡ��
��:>�63����ys�����0qz����L�Q����Su��Tq��~/�٢a�@U(�z`�Q�-V���'�+�;1�R^�u��I���~&FR�'�0.��[w�6�W������
�H���nq�dL�IGhf��&�,�%@��$,���h��Aʂn������e��3�����d�|D�(�܅�,���$�""�oSo��������!҂9^��A�V��J�;n�\[�G5�܉��l9+�w����hr�vHLf��O-��8�
l�_>��d��e���*��n\p���}��pȈ�$Fj]+�)ww���f����� �<_����6qƌ+��ZS�TR P���hS��Ϭ�l����IA��c!6�s�"`�1N�:�	ntĴ��S�o������h��� ����5�76�O��8��v	�*�&�VEY���R֪F��glt�KVW*�����Ӱ&&0����و>�{�q3re�1�yA���A�޸�O���C)n���7fo�FL0�x<t�%7�.#q�K���C�CC
�*��LR/ r	s9�r�{}}�l�-d~^4�<�ӅVx�Қ���e�fmN������QCyq&����b�-c���cr�֑�-��(���8�
�b����������e�͍���'��d���wY���Ap/�=�:��Sjz�ua�t��=��ԕ5a�Y��I��N��,���D47��Ex铙:> �0 �� j*����U�\پG�TӤ�V���=�$ɬ[7s � � �U���Ӗ��p���aF��.\E�nE�ZF�v��31.rb�L�U�˕v��2��]�{l�8� F��nj͌6y#�}�wJ�|2����֏*
�J:�L��óB��=$��\�VHP����=�d��pQ4���a�Aa�.1����_�7Dm��9�&Tku\ ���
��A6�Mh֝��+�b�o����"�p㉜</QX�(l������}�UF�<�ɣs������Z`�\�@��u�hJW��D�F��b$7�'��H���c�X[Vۛ[�q�!Qv���jd6��-��W�"����	P�
'M@�4w���*%������'D!�.���������/+b�Z�y$<�	�sWFR�����4�&�&5G0�*IN�}F�,Ӛ���!�Q��n�2���ծ(��a��/��l��#*�ƛi�yh �<
di����pn�et�`+���3r4�cK���5ꢒ��v�`� ���,{��'��،��p�*�Z�B.�����Lgn����J�j�j95ˉ7��_rH�@Np?4��K�i�J�4���ȝ1�"����].��r>Ζ�	+��%,��w͠+f�2Q�9b�d���P8�Ep����ѐ�B��(�#�Z-Bk���5�%_��O�$lc��>�Q�4Pj?!���i��rE��M���*#8��m;s:#�����54&H�y:N����TszrPS��u�ٳ0_~קWZ�cy`Uf�>=��o�����=P2��ŧ�x�V�+x��A����x�
-�Vi*�4�ź��"�5���� �j���qا�r��֌��e˂F��)��� -��*���:>�?�{��O&,���r��Z()]� �U�/j=��]K��k���t)��-�S`��H��C�@f�T��l�]��PW�&+��/��x��f�UYX,�V]�����M!��j�������Z�h��jɢXs�X��b3D/��W,r�͆0�|�R[���d~PL��Q�Rz&K)�<b��>�E��'QE�'૛����s�HS~�mna���@%��xz0��4��W�f�%�9�zS�ڥ=�ia;�H��:���3z6�������i�n5o����A!��jǛܲz��{�9)Y��k2(��w&�;�9����!;9��H���� ��2����a"��5�g�.^����r��s�nk�R�V��1�
�2!��u���銖����cd6���+�ۅ����)�lˠ�ɠ�Ppl��w�d��d�4�bD�=��C/vl�-���T0�<�bD-{�R]���p��F��|����V(
�3Q�B9V�3��T�:{��:߁/��,	��xlf`ݎ�R4����~�a��A�����?26��4V�o̮a�s�&��ҒAo�r��7�v���]��t��Uah��s��)���=}�-�S��2^#��*�~�� S
�yϑ���/i9�wU�0_
?�{�+|���R%��N�{ IsT������Q�E�eM�c������4&���l��:g�[�����.������+�t��(w������4�*�X���@'}���j���'y��
V�M]��I�n���'��r�J{����d��Ŵ�v���%H�d�]c\���p���F%�RyT�2�8�Խ�����ZS���hba�W�-�:I����Y��$�ز��lNf7�gD�5��R�P�g���(Ŏ��~/<��FGD���e�>��������]ņTӂ,?&��dH�jL����	&�����L5��G;/~���8�aQ�͆��u���f��4�{o�V8�sgV� ^��!��*t$�0L	�����;i|��(:/O�/:�~�M���3;1�?����ul����^��%��Yj Oeۀ�P�bA�����í%kU�����jk]�>�o��)��I�6Es�
ki�{�f#����I��!/�C�3R©�E���f�t�M�����)�����VS��j�ut�O��|�;�����<��y�q�)����:�{�K��	�V'�ńLԡ�����?��j^��BfV�Q��&����V�@L$i�|�j�j��RX�b��a+� ��k�Ҿ�Ý�EKŋPo)�=i4�0-ʳ����i�s������DA����J	S�*D�r�YrG����ZNR�M�L`.j�� &f C�nf��>��w���:h�qd�Ϫ݌)�ZB#�9xw��K�UM1�֊��@�`[�X8�bE��m4�z:��}���mP��>;�;P�|):6H&����8'�����oZ�n�;6�H*�Bi��� $W2��A���\� (!ε��A������>)�.�,���A��DN�Aw��@�j<K:��M�`�(@�=��$0f�D9Ԡ��@w+x y�|J���5�����{�?�'ř�r�}�bW�@�*�g�B�a��6{?K��E������v�!*�f�0�)���	8�����V�t���ɻL�vo�J�R�uc #���A�mĊ�x�	t�*\�-ŵf���S�=��x��|U�jm�=��X�8�Tjx����ZdYX���֩DxCJ`�����q6���B���M��H��a`�YD���1@�C��%R�_C�z�b=>��qT�����?��&���ܢ��sU�,�J�;?%� ҎJ�}�B��`*W�Tܲa]��r����dRN��B�i��hC����#�
ف|��qܬ0Z���P<'9����i^�j&�D�Ͼ���0��F��A��B\)W�]5#��!���ƌS	FB��-��?�ٵ���SGp�Ñ�	xNp�Vl_�;�W�QM�ZltB.�A%r]t�G��t��:����N�w��7b:Y����U&hG��E����Ӆ�⾣ď��O$�X��5q1��)���b~Ov�Q��>m����@V��V9WH���Ε@�a���$3��-�v�SkM6"������ � �{�ܒw���6�XS��EH����U󩁜����	J)�mq�1�P�~Ll�m�1����	�&�K�^�q/�NBcX�R,=�p��!��H�zTXp�EL�Q�9�V���\Z��+]�~g��.���:?���%7�O�'�5��R�f��� Ă�M�(�1���},���=�ck^�4P>�C�I_)��O���#�q�d��űiX�D��EW�P��+����Lq͢> �b�����xj8��Vå�+�G��������/����!n�φ���&��GR�=���=\W�g4��a�?��1b�1�\��j����%��������3-��m����NG���9����?Z�̝zAa��^���n+�ۆ���7���]i�#���0&&f!�1u��{49=8�b18���L^#��?�0�i�3��=� �{=Ѱ�}���Eb[�	@gw��8�hqh��V5Y�������]�*�1������7�Q	6ɣv��Y�����E}�3m�c�~� �`X�L�s����_�Z1֜[.��&x<����M�p�k	%��O*���n�h1��S� ��3�a��8���?P�G����Q�����;�)���zEI��;��rw��Owȉ�azA���8�=��]�c�&�ga�J����Q�=z���?x���$�4�u����t�d�����?����pu�G"I�a�M7E7��'zQ��̅��i�J(������5l��{O��H�K=��(���d-@������"q��S���1��k� �3�$��b��+�`*oO��a�i.��i.��'/dĲ,�-;K��nna��4z���3Qm�ʄ:#�d4?+9:Ve�S��A(�B�Έy��c�b;� #�A�{�Y�zC��L;�K��]�t��0}�7�-m�v$�����S���N_�e��2��?c}��H�W��� �A@ėW�A�U�y�W]�_��2V�#+����5���`%��J��p����E��</"����1�_(��Ѕ�W���0{���g�䘕I���0$�����Q��ə�͈͟54�~�v��Ԫ�򫛳��h�r��WDٝb8��`�ܔi�@��������q{:��e|� h9c�[ ����~BC^ϼ��Q"��i�=��e��Uj��v��x#�GY@���tS�&�'l�&ʻ��L1Z�nd��W�R���k]�W�GL�7�����s�>�SA��I]m�-����r�B3��4��'#����{%N]��/��f�6\� qO/��Av�L)z8<e@���~5���Xi*�
n�rwwY�^�ߨ�2�t
�-}�7�3H�]u��Ķ.����=f%I�*N�c��3H)���8�@>�`��qu�mV��xz8N���3+�_g�Al����\2Bᷩ؟�\����1T�$Q��G	�y~�c��6b
%�=�n�h�����"���������ݬ�-h����_7�n��]36-O���Hq��O�,bE8_�:��^x���	�GPO�1�B�&���H�y�=�!k���}�^��p�W�x
��ҋ,x���E\ģ�bYIU��!�c�-�b;u����o��3I3!�|��ݗ�~� ����E�[J_8��(S����V�B�
}���f0"�<ĳ@�*-�N�e%�MMKr �M��7��#�o��-?�0
�&e�y�bgEH��ay��I�1�]���$Zy��d�b�-z�M��c��~SKfv�t��c���ޖT�H`�u#�6tY<S����VA�߃�L���%���ǥ��
�,-�rg�����eܨ܌cɃ�jX]�m{a�[�J��,8�ڮŜJ5�u���&��+�5dSR`���g��|�wPrMv"V�q/
�0���C6U�ܖ��^�~]��/~l>s� jY5ё�6Y+�k5���������Ov�>}�zI�Iv� ��w/�r��¹�6\Qp/�&�OiFA>��z�{���~�|8��@�F��
,o��M����(�A���߲a���fC�����{�?�	�Lg����.^�;�掛���$)WÃۚ-9n�/��G�I{�p�3|��E��SԲ�& /��a�Q�ضc���<NZ�djx�����c��<�5�(����{ζO��R
�8#�P�жEaQ�-c�F�H�����X�X'��	�� �� ��c��C_�#���'w"����]~��f� q�o|����@z��Vފ���]��C�xq���2Ft�R�s>�_(O0���Λ-j�2)���O�"<Zq2@�\��E��z�S� o��-�VTcͿ�SN^Z��-�2z����������C�/1�Uϴ۰��$�ղJ��w6�%� ���<p�N�e�+`��>:H"��0��&(RF:#��~���,�������r��NV��Q���M8��`jQ��g������]��Ey34�yg͏��I�7�h��?�4n1���\��@�[��P���s�^q"J��l?���vfÌjYƁ8|sQC��ԧ�����Ik�yd���"��\��a��Ue��V� �u���Gb3��lR5�)×g.�-��Pލ����y���ۏ�ҫ��� �q6�a�ح���B1�[�!������S���hVi��o<ߛ�3�i�=�y���K�-0�X�I�9w
-����d�w��H�B�J�Վ�b��n�XH{7hw��MW��C�I��������"Lwgh��jrW�v(2��O�q��UW�;�\^�0��LcW��źp�&��K"zK��`�,Nm�EDt�o�Q�^�6�b�ۿ��5�h��{��2�ަ�MS�@�k�D�O��Zi'�3=�Nk�YN�����_3lN;�����M�'���b��o�_8��qT�y<)�ҵ��Ѡ�2*K*�J=C������/ނG$q�����?�?���U���"�P'_\H�U���|�Q"/�ʖ���Y@Y��R�����p19u�����V-�\RN�>����9s6׀
;N�����^ņ*t�AaW�F�z���M�D�
�KXS-"zD\\���YSw`u1�0z���Ֆ�z}M>�9C T�M�]�y?u�yl�?�CT5���t�����H��g�uM���?+�:�u�N�����[�βT��,�òy���Ƌ)~5(���M���^�ˎK�;R3�/�7^wW�zH3�]�I���3&`=Id�L_�}\5�ڄ��҈��uy$T��B҉>��n��里ދ��ƢY.+w����zht��j��PާI_p��R���0����vGD��A�0w�L��7o*�eHR��O����&���L��j�%�Ʌ��Ιz��s�� �ta���{HF��Cb+ד� ��_�Ksq��^~�:'w�ڊ���8o̆����s� �+G\�cT�XU��C6ցc��-GHEº�aM�zR[}Z�?��-jA�X����?��pz&��������n�.�*�͡4}�1�ņ� p���%��?�mt�DG�j;�W���2:�hbw��"�u�%P�-�6���*Y��f���[U)T�����N9�!߰������oqG�j�Q��23�����k�]"�mRv����Wݶ}bj����0�Z�LF2�.W�-�CM�GԤ*4��W�"H�ўa����؁s�׽�bÅk�N�t<m����?��k\�2��'�ֈ��s}Xka?�bcj���0+g���A~]�_<ca�]�������L�+m��"�*o&b�[:HV�pI���}^2��h�������:%O��-�����]�ш�i�@���kқP�8MuD\�K�P�bz�����1��
M W�^��	ޤ�Y�� 	<��'F��q������o>hG�ۅ �`�}kO�+���q�6�cG�Ǘњ�"B�1��*��X&Ƥldo���h�ѡl�@XۘZ]&U��QHVa[���ׂ�U���ZMC��7M/N&Dۭ'4iN[S�����\59�c�Q�3E��K��z�&CV[ ��Jv�@�E|1���D������s������%m��<�~M����� �����]p>�|�v4�pQ�L�+��f�hHP�)^:�:yq��^�,�e�vo�F�ʒ^CԐc}�->�IѦh~� ��U�Y���s;�32�bS!۫N�N�5���:r���c*X	S�
��3Fr]���ȿv�on*� &���w�;�W�ZC���Q��+jrZ9.��l� \��Q��o�_�3�gxwp-��ҭM�A�2ف���>�F�4���ʦ�&�AGV�)� 4�6o��r3�%y�y�4F��$�C�S��AB�����U�ҽ�b"��#|��Đ\���>�;x��`���"������qD���fV��E*9�C��吁낄��j�����4m�2f�+������}?�S�'[8m��u��=��\!q��ZX�'�������0��Q1�}U�ND����XR��c9��>'����\�	��򯤺�2�/�}�EZ
��L��h>i�ھ�d���:�����Đx7�8� �@a��Y}!JR��~�)��}�j��]�(3S����}�`2e���R"Sm�q/�
�ﻈ���Y?J	Zj�f�V���t"��"C��	�t��BbU�?�ʸ���cs%q3��13��̇���q7��|�3�3�|A��_Ԗ�cԽ�2�
��6k�5.XF-�(xn���l�
@�^��U��?�x�5Q��<��9q>�k2���>�˶���$�@�(�g���E��̲���X��dn�����:+>d��+��Y=iF�QH)H�1��nD8y�u9��qMˍ��#�H���݀@�\��t��ؕ�֪ID5~]�\����a���0��9x�����Ёw�</��p,8|�Y�̥��u>�1y�����K�7 �n������L=`^?��s��B
M�0�Q�������=�0���c�ʚ�8)��Ϙϫɷ�e���Gx�`���+J�dS'��(/�����mڛ��ĹJ�]�n4�1���<�sQ�0���"�e��z���+챦c������4;�mȉ�mv_��J���ˀޗZ��Q�x��3�N�}�9Iu��ʴ��^�Ȱ�b�������D ���*�%�p�����7��Z���WYB�䏃� ��c�6Wrw����eR�������ĞX�o��^	Z4r��h���]�tua��9��_��_�z�ܛ��RX��U'�������=����$����y��l(�8�A�\�;qږpö�]r�o-!ǋ~9�E��;�4(#��sr�F���+�8Ē�b%����	R��̻Sm
�ŉ�	3+�ى�跔G�M�0 ��J���X��ZZ����݋D�˖���}�����+Rq�ِW�
��;@0wBa�Zb9�g���h@��]�N�i��u�F:�/QbGp�K^�ǚ��~Pw��;�!Tl�����t�lx���6cv����f/��F��B��Ym \�	�s��,Ɍ��^'TK�\��0��D����Ƚ��/z�F���C����CdU�3y��.�+�>Z�=��y*�G3��SZ�A���27�6a���,���G�*���7���|���d.��F��/_%w)���;���t�5zȭ�b71C�I��YBW�q��ábg�YQ�A,35�s~�<Z�a;��ݨ��U��qNױ�WB��uekKyiS5��� �t����v#�mSp���G���6
$�1�)�+����r	��Md$��,5�����-9�+�1�O
:�^�i��H���$*R��E�XȤ�{�g�f�0O&���E�p�C�X�3�#�<��/́��e������R�ҝ3g�O�gv�j�~9��FT�+D�4Ir�~a����^� �1\vEnQa���hW���2��5F�f����B����1^?
�r(�V"
b%�֨�m�!�Îf\*OZu��y�z|*䪢�2bjO܍"�h��Q���|�ho��`��e�
��ȏ(�Sܚ��b���ZP_�?�z����(�Kg�.�h�3���ݦ��6�C��8�?}<���O��b�P��]?�ol�����rbE�[� � ����rH�{H7jQ%]���k�@�����hn�u�8��W���R*~�4�8o�7>q�U9p<n���ԅK���v�(zr�4ur:9U�
��8})�jJs���}��Ā�o�
���4� 1�['�q��6AN�G��(B�!v����`ތ��vos��Q�I �~> �}�g&_�0���`��#ѩ���� 6�IV�����a&+ϥ*��8p��A��o5�HNA;��TQ���!�� ���%I�G�!��"/iX9f�)h��{h��m������N,V^�tMg�R'R/X����o�wF#p�:�ߙ��j/�;�T*�m�G�� �N9�Nj讦�s�6#T.F���'/��k˫�6���jx [�FR	.v�D�!;"��@�N6*6�D�������J�:�����NK�rkH%�9�����deq .��#�YMp��V�)�M��%�U	;Dp���O���q9
����0+(������z�b��̰KL����;�g'Ѭ�~���c���V�p`�i�`>����.��WT�:�������5���MӜ: ��Y��Q*�'Ex������;�Mso���
��)�Hi����W�s���
�,c6��|���<%��@���ҁ���1�8#��:�&+}Q��eS3�*n~�7ր'��=%��k}o\�1��n� �̒WO,����2}�&������f��R$��(B5�����hn������P�6\���o!�Z%w��b�V�)�dFl��s����g��4��ͥ+v>@|�t6Zz���W����<���'�����
�0g�-o�GFrK����a����i��b���U�&���jw.hhX�"L2�%W{����d_�%��Ev|B�V�iyh'Z)则��T%��E��.��c�?� �W�LT��Q���sV5��V����|'ҳ�M�:��K3}^g%�<8~(. )9�$��<꿿Su�k�qh�&uK��[�*V��d?�ɭ�d2�L�[I��]<Z?ֆ�Vީ�Ck��/wE�40a�Ɇn����͟�T�dk��P�S��s`���!(����:��ҝ3��W�ń�q)­81L���0̏����^�M�]wkV��r+�m�t'b ��/Ŏ�7M�-}^\!�"�;UZ���,����O
��z]��艭���7��5��c�ӣX� ���Mѿ/u�.j��R�#�?ݯ�K_ң�KV�c���eZ��	��|���A^�'�C�ca�5��T�ڷi���y�����>2�,
dʹ��ud��T��$U�`*�����ݩ����|6c[��C@]ε�B���>�AH.��-�.��^ R}nb)a.�k���ݓA�x�f���w�	����s��c3��� A<3yN;V�OV�@}<p<rI��m�FWu�_�0	Un��w�e�^N>цf�vT�Gga����+��c�.Vp����h���w�dm��[�������ʄo�~Pٿ��=����%��C���EW�Y"@#�p��O�N�g8D�b��`b�e��'���̘3�bnu�Q+]��S��ŝ������qNך�r���BH�L���c4-���.�g9
�!9n�t�%;W�S�M�T�q�K+9?l�����V�֟ �2H�&Tl���2u���S>�y��e.r6�9S3]CB

�;l���p࣎C5�����w9�*������A���� ���篕=�6Ұ)_�[`���O��FE�����*�[���U8��<�� p�Ow�U��#u���/5$ ���b�n�d�S�}���.Z����`,�;��i]���n�Dϐ���^'x|��~ߪ���u�_�!�>�S *�9e�����GY!��Y=.���]bW,n�e�vN����W����<ֿ�2�[G�U~�Zc�^"�!���Ҋ�jn�3�{��������!ɸ�SO9�uj)������k���$S�޳�>��m�ޡ�пH���]8P����L�cQP ��!ß��g���!Яd�kQ��Bd���L������]�<��af>���o��Hp��}g�t�^5����\�e��2�ʈ���Q�6�ߠ��|��ج#w�>��px==����[�� ��b\R8�(�p���O��b(U�Qu�A��?�<K9=8肕6��ݘ�8�iy�n��T����t�ڢx�b"s���J3��3փ�f۶����V���7�,k��i�{���D8�hkx���uG2`(�=O�^P�9	?�)ː��u��BؤA�4a���%X^� 9ꄋ�������[J 2[�s�� �A�-�-�z�Ն��673�n}�t�BA�Q�r��KYx��1Ȣ���X�y�u9Nu��3�\�������M���X/��c��=�@�eI�,�)0��-@�!v��<?���g�},�-��f
�1�"�sG�6�� 6��`e�Y����~��p�g$9���*)<���$�q�Y�EA����ܻJ��.R�GL}ij*�P��0W��ࢧ>����@��p�o�^��[ڐ�F��@L���)���j$��v��d�n�~3Z�=��h�r?��;Ul.vۦ��?�G�\e?B���M����]�eøM ������%~|�ߙ�u90%��Jd��R�XkA��a�摅�}}E������m)ex���Ⱥ�I$~cc���
��o��85x�\{';�v��G���Q��n��z'*���Z�LT�n�ҒE=ݸ���ؠOzJN6b�~�&T�Y�7O��峦J�w�rޣ$���b�k�ES��dȘ)<��)�s�grs�	����݅&Щ��;�o����L���1(�}v�rnz'�TN�9���ȑ�K*Hd�|]]A�=M ��CL
r!<���W��u���:�m9\�ʟ�����?�<Jן)vψ�8��&�/`��9j�kq�^IO��~�%HwM�P�#u_�J4)��o} ��0���mrݿfa�k�B��1��P�<��f��D[��%w��g�ք���NF����o�\��G�3	�F
t�K&2˹��i8�U��BJ��������V�6�y˥H��XEn'+�,
�~��y���h��g�W�v��3����u�S6�wd�����4��`�f=�<�c>Ƿ!E�>B/}B����5[#���C������=����߱��v\��ॴ�~�:Y{Ϭ�H��0_�c/�P��  t�7��*��J�0`A���T�:n�7^�O����1l�P�6P�3f�����`���S��������iCm��A�-^�9:�������j�{��p�U~} '6^Bp��ZZ����%Hnf�"��ē(B�r���J���9��ꖤ����:[*�N)`q���#��x
Y(�p����W�j�^�a/��3^@��挸\�U����L6�אx	��	�B�R���f����SVz�<�/-#��?��jb[��a�����r���V�ba>�iW������C��hy޿�W�A=�p-s~Y��0Q�gN�
	B��áx%����5�	�f�n^2~�f5C^-�ͅUH��<�g��j�5�I����	�>�����|����i&H^f��S��r�$�fj�5T��#F${�R�hY�.eYXI��Q@��.W%TM��p��tτS�� >��|���ռ2�ηw�\W��'�@���2 ^i��YskW���vI�ƾ<��vh�h�?ʏv*�2�:�@tD���S^rۑ���O0�:��%�	{������oOƒ�G:�L��tO�a�*td��V�����NV�*���Nh���WlH�B���~�O"��;�/��R�8�
��ڝqq5���=��2��D�c�hF˷�����U߉��������4�ϛg��k��DC�`ZdJ:��2�m�!ײ�z��L��k5�eP	S-̠�ņ �m���������ֵ��A�y{iR����}����`t堑��v�e� ���+�����>crT�}��D��a��Q��J-�sE�S��ʎ3ӳ��fg	/]��MQ�&Ev�E����ա��-h[a��;Aby�\�jB�害�>�z���Q�� �s���9X��}NZ��rRhK�����|bw��`q�r̽(�{�='���{L�}��@��g�4�[	��=[A��h�-h����?A��� �@�`rJ6���t������Ze5u��^-������6K�%�����/����x�^0��a��W�����_���-�:J�lG'�9�
A0��2�<51��=��YԜ*�.-���{F!9R��[����1�$T�$G�%l��Z�p٭a�X	�oR���q|GiЪ���_`��Y�G�lT$V2IܘYll�0��=� �g�|���,Z�!sd��18�N�gy���]����<Kz�`�7mзGW��ꂉ?b�l�L���P��5�?��Ni�e���%{$ʍ�_j��R�䮉�z�k������ߛ�`�Lr�3=���56G��z_�l?*�y��{.�h�����|�z]em�g*ǣ/'���֩��r��k�<�����i��e����'�b�$��+Uh�j��C:��R����de��IX�r�Q���F�5����B�M��Ϊk3a����:`��o��$Q��X4]����;�X�ػ7����+pHu�J�q�����s��#�����_��t�n��ae�+�k�DEf}Է@�Cbo��?���j��������D���˕����/�}�EM��en��sqD�����54=����t���0���E�5�M���_>rM^�n�@��߬KYh#���{�ٺ��"�x���ND���u�#��tpCO�Q灭N�Fbz3j�ށ�]}2�"�-Iz)C%��[���?����M�fu�&�3���:։ڒ���_��?<�"�l����ʸ�iHȏg*5���W�{T��.������:�e��:x‧�m��DO��fI� �
��T�ݘ�N`�ˠ ;~�N�ƙ~ڦ�dv�D�� �*���NƩ��ʬ��*V!�&��r�8��v(�i}�6z>�@�F-�coQ���b�4ִ8����i\s������Ι� #(�f���U��b]n�}{̐o�,���[����4�Ls�U�nm�@q�LT�@Sx U�	Ũ3T��
s�Dw��l�uoĒ���o��A��9gk��VAw��z������cM�~)��Hپx��bKG�m��,��rs�)�i�{E8�(t���~A/n��IQe�R�^ġg�	gk�i�6��S��~,;a����_֯/N6m��׷�Y�dZh+:Ug����X�P�[��E$.ϵ�������`��8��Q����*��SF��o���q/H�8� ݹw`/��<�� BV�6$��ڃ�F;�yl�>a�:�@q�gj�{'ٕRWEu�K��	�~�R�46��Ɲ.��A#B�������C�3��g[�,���x3����J��?Uw4����XQf.v�|.��WVY�#?����|��@��M�Mϟ�z�}�n�����8�HGz1�J(�Eq�U�
8���=o���D`�lw��^�nT$ebAu.t:�G���u�sJ��+t<y��y��݆	�*�ʠ�\'�x����PQXֹ̢m�@��v[��f�yd��S�W]�!��-�!�UI��8bB`]y���v~a|M�%���z�52�8��z��Tp��ihܔ����ǰ�9-ݑ�Rig���.�r�a��o��
�ђ�Mn|������ȳR�� z���²W�;IgoA��&CF�� Dv8/ �q������jK*�jY��F����^��3�^�D�vN��b- Mһ�c�&��M7�Jc_,<*�\��C��P��y�;b⹍�"�H��۰�b��@�<:��8,��6F�	ޛ��w[�Fn������)Q�/�@���зJ��I)u_V�Qs���HwǙ脏^�\l�����%>�{�ae�W���S:F�{�G���\�� ̜E\�&�HG�P�gd!�X)�����B������y̸U�%�9ho�c�,��ur\F7/8�"a5k8h��{���p7��y������<+VOyF��6���a|�5RRͲa��?��Xk�PӥڋW�m4�:&MD�'"���&s^!Q��8!�KI���: �;����W�zg1�"���>���Q����0:c���A�T�H��TD=�p�\���3��7��9�.�҃a�	�r.u� (��<���	�o�����"��&��e>�$�0�o�X�̀��de����`6U��J�
hpx�44M���#�h#!�ڍK���+vo
/Ҟ&)��}rJj4�9�PU��\`]���\�g�ƶ��䪴%9����,&y-��#b��/ቮw��e�Kjc����
�
;$�.�R���-xX�ogdDv�Hj���:i̘�j��Q�I=���'|��K�>���
\k�Q%AD�n٠&�%�J�yZ�ʑ���>foy�dAa���t��r�?v�@nmc��v1^d��^�p��AE��%}�	��0[N�dܮ k�e������\r��oI� %��/I4��?��x���C�gp!���_1�� s�H]�d��)�m&�pi��J�5��`�_ �DEF���(R<d��#���	�yX��'j�­�b�(>>�
�U�i��y5�)!��FC�㰆ͺ�K�L�.� e���9�V$}dvy	��)-��掽"�<c�2s������z�E�:�j0�o9��G�P��G׷�]��vk�f�U�{�&rH$�D�L8Y�Mޖ!� ^d�.��o�5,Y���	�{��9�M�.-���V��4�>�*�jB��%q)|L�m��H���^��/evؐ׽�ZPu�����/C���5� Ş�����f��,U׃m��\���YM{Z�p'�����VS0�BN���Eb���;
��dg� `x٦&qwc��*p5�����K=�b��[�[��RN۞��T�c�-�ܤ~���e��U�	�[�b��_Qw�5�m[���,7���v7y�L�J�a��n����ܽ�[%�D���h�X��o2ZLN-�H��,�	i�1��p�{��f��gn��'�fL�#2
Όr`=�K����
t�����ꑖ�������2]8����[�K��Ԇ�3fI���'\��(2V咢ik�X��"��}9)��,�?��/�K���Є���`9������~��h]�^�2��V���݊��s=,�y0�/�����l��B�a-�>J��|���o��j�� ��O��P|�\i��t�*1�\[�d�)������>�h���»����ށqZcpn�Uˀ���9�潀�$ & KŒ\�}�<�����X�~>�*�=��s�	F���Z�� ��Uof9�r%3���l�����%np  /�@�e�j�~��N���
7_qF	�%*'���*��R�T�9>,A�ׄ6�	�zb9�o?.݆`ݱ,_���3}f�P9c*m�E�d�O��k�@�ŤM7G�)/L�;'?Q�s�'�y�`�ⱅ_�g>Q�b	��c;��m���]ך�d���b ���w��]��9��~3^E�">�qJ2�)�`X&eW��$���3�A�:4�A\�Y �x��W]�Fd��g�Q���P2Q�!�>���(��^�j����?& � җc����Ū͆a��Z�Ĺ�[Vw"��ɰO<�2`���?#���/���֮�UC�.�8��2�>֌}���bzOq�Uhm��j$��&�r��f�"[�B�����Q�����f����ơ�J��������#9h��Mm4��+�&{�1(\8��q!.�/�X�+.��k�?;�t��Ư/fi��
�.��})H/�!�A�4a��X��3a:kC��6����;���e�j��D?�:20����L^�"��!n	��L�x,�Bu�#�x�p��i�dQ`�}�k�.@rw㫋l����
7�T��.$��L�Gxo�L��kƎ�"�lc=Wl���-���#��a��?)�&N�����,���*�Ҝ��������S��O}ĳtΓ������"��i���!5�h��!Ϣ�?I�9fE�#�5w�{�姱--�?�bALa�x�?D�!I� 
�,�u���҄$�g�撹���Uu�X�K�\&�����'��`K=Psܧ/���
��D���L�Ѽ,���]Hf�O���q$�gƬq����ģ/�$,���/�ގ�l�ַ3���L�	e�nCӦ�;Hɱ`�L��4]ɲ�ʇbt��J� �X�W��f�n��(�0W��Ycf�$/񃍢��el�~��Vw?��׀Su��,{���1�����o~d��Q�9sz�!�<�7���,����~�X�J�D��������
��nU\*sp��~*��Ki��B���W��~����LMjD���ʳH~�aG��D���i�ӽ���9@��`9��G^��a��3;W�>��ZZ�0`Ň�u�ȍZ?�{��U}A7|Lu͠T���.
_ՠx�-vM'֮�PBj���e��@z�_���\�j���!�:&���2<-�%{�h�V��L6&�E�[SX���5k|d;ta�0KߊD0m��I��ެ�߹Q�s�G�IFl���m�;�Zٟ��3vX:��{Si� F���
��vER�����ec�V�׈عU38+�uJ�D���u���D�L�\��`P��|p��N&Kٚ�|wg�/ϼw�����$"vԺ�I~���YVf�_��V�>{c�K�H,�k��X�p2�V_AK�	�ıDbS��rIt[�ȳ$�f8��rFA�Q�F��[? �y�`���M��=B��Cq;�a ��o_����7��y�j����r��}-�a�0*���`�/�R�����CO�����)B���{;bX���B)�v�Z��+r�s���:����Fb�Ơ�_q�t��Y������v��3�$��|��3.qTS6�"������}�gd��%�-��p��ʣ� O���ҤId'���LIP~$C���4���p	����V����pm^��Y�{��$u}H�<���G�B�)m>oi�,�6SŔ!S뫷�<�ؖ t�i�
u��fWƇ�eZK�)�&x_(�j�ʋ����2�W�
�}a����+���W��-'����g� �����en��ƴ�B�)�\ 3�6�O����M�S�N?�D�;�֚�=�h5�Q��|��cZ&~7�ma	���E�p^�N��� ��9��9��'v��s[բmkߝ���6�S���A����$DRi��X�ռ`���[b���q]j���ʳ��~��8��c_f�����aِQ�m5E�I/0I2��如�Y|�V6nѐ푖���h5B�C#��ڨ�+�4ٴC���{b�҃͢�.&
�3pVb�q�y�By5@C'{����Bܿ���U��>3$}�xB�H�7h���[��9,�����>6������N�=ӆQ��=3��4�!� �p��)�E���-7���x��1��#a��P蟨��Uh�GB2
Ѕ}e莉v��vCA3�H��D gl�e&O�u�Pb��!Gedɭ��'�9��_�s̰ڱ��NRgP�{^&����U�R��c#m' ��tx��i�6+@�态2�b�,è��j����qm	�lJ=�,caW̜�����\ոW���Qy�v<�J�Q�����H��0����ݴ��g�:�}5`!�5�6@�eMO��/t���6z^��>Dy��H��	�[�Nl�|#�:�d8z����u�Y�r�d�� ɋ.!����w��-��d*���ý�ȕ�.�CD�J��3�B���k'�9�hR�����������3Z����֫C�]7���[�@!�3~����N�+��]"%�ؓ�F�4-)dk�����Wn�/�;B��>�L�$n�e�����o�(�y�f�d��s��v���XN��`�����
-�"
R:���[D�+��E�˖~nۺ��D����DT��9k�?�����h����>��F#Ш�濆	��s�� ��>aT1��U��fp��.� ��
.p�8�-@��gںo�2Sm����.���h��O�y�
���"�\�Ns��<E6j_�.�]�I"*2+��`)�SR�����qn���Q�7f�����L�i�?j<m�!i2e�ԕn�0#w���!5Z�ɲ>��ե�Cu�_�6��&i{3q�eb��Z���f��YWa��g��f�A0�1��Ma�ף��n"��B�ă`���\(�|�(��I�~�ʫ�&�m�u�LW����D����Y���dy�Q���6(���(��R�;f�f�p��y,lH�i?��y��w$�7J�b#'�,�r��{ٓ�I7�?X�߸77�l��\m�<�v��Kb}~����d/Z�W|��7C��@ݠ� ��ɂm����Gwy^����#YJ��8g}B<��&k�1z���� ���ӟp��D�4��9�ND�0q킹1�vk}_t�a�(Uw���9�)`�x������0o�|- =�ʾ0���b�Y�L.����y��=��9�	݋�Rt8�_"1���QMs�os
	�E���.����@�#{#|���D��cYƆ�y�{��7�뜣��F����b���[�>��G%w�(�?�1k ��:l%�S������9���~F1:�H]Y���8x"�1���ȝTv�"t
4�e����r�d<֫7ˆo�1�䌻�sN��wR��<MSu��,�\��p�*�Kc{@鵵O;�K���=�*o1i����`��8ߚUX��9#�6��˲�(���_��+xm���
|�ߝ�I�4i �Oo�	2o�y
��}?���q�J{��Ȏ�7��ߞW��S}{Ev:�ԬT6���(��-����FeM�]iǪO��kT�\�㥥�N3�ǔI���;i�;�8�M"�	�Af�V�cI�]u){	�/�v���oįV�4"�~%��	�Y􉧻B�<N$O�I&7䒼�Td �~(�b�5�gg�r�$1i^"�Ƹ�o��:P���
���%x��ЪP�ۥl�v�8Cvܟo�DM�����X�H�T΅�7t.��qg�)B���É�Yހ��ْw�o�����p�PK��{�o���	,�7�q��
��CgI��8A}�B��H\���ZKE�+ �K�c���@i�1X'̞�^T��3lt#���QQ�s�%������f3��>�\�b8UVx�a�?q�T�
�����5^F��j�O��9�?�g��K+����x]Հ��a�(60׊���M����a�N3{���1,���'#�2?�=?�x��bb���"��vB���)!�U��~�]tNe���\�ѹ�G?E���S�|��tB��)�"�%nѭ@:%>��&�9�v�
P����d?BV��X�y.�(Ԇ����ds }��&[��g��NfC/�[9P8^�~�tij�a�/��N"�J���jd��SM=ŗ�|��Vʎ�u���� �Ƨ�$i �/�>��D*��k�Eh��0��<����0xb ������עi!51�@9+]���s��B��i�/>���KduF
$��E��1|WK3����n��U؎6Ae����s�M�B����LX���fApUc���[Y�����}>t��m�yj[ PqY&Ei��11�9(�Ft��CP��V;:�A��m+�z�Gٌ��O1_,a�E�3�g��x��.�CxDqBk�&k"�w����u���˥o�@���لoëv��v��K�)����~[֌$�t���L�'���HQ֝al�~ω��,	/�69�,7�o���ٲ������!��;���R+g�|��˧9b���4�Kk�	0�"u�1S�|���]2�osb�"������]{<����J���TUE���e�N��m�!]E�Վ���y�Kvj��)Ƅ�H���[d8iV$�����E��������I�p�g�Q�Qe�6�m&mP_�r��C"6:Z���})?\P�C�m���}ߐ�a�s�J6C~ a�̵�q#[��۪�@�ȉ���HM��ڭ����ʯ�5ǕC�ujM�xK8yܭ4�4�J)6뽒{�lJ�8�]�ٺ�4 K����ۃqFf�ٷ�o����f ��eD�»��oS6Kq���l�o3x��]���hm���e�ʌu/���e{�˼�Uq�(z��f����ܻ��<��t��7e�2�F�ō��y/�,����G�K��w��f� D�
����Bt ��� _�:�T�[`>h�C(n_�l{v��b�?�1M	�vQ�8�줊>����\R����$�u�J6K��<���8�H���E(����*0�����~���(4��Fg�v��J��[)��~`��E�Gyv8�{l�?g?Ϩtn���}=��Tb�g���K>G�m�Z�	�hoU"��£
n@|0f�)ț��9%
�S
)]`�I=�A0_�Q׀r�k�W�P�J�V�H��� �:F��!�!0��pOr�%�G����u�=����B=��Hs�<m�r����,��p.5l��ε�h����T��g���T�#�M�X7g� �_O��S�́�hj��Ǣ�V�����9k��p��ͺ(  ��Y@�����wɕ�&���d�n�z�b*�����EsY�j�*ACN3�`�|�ڥYΗ��vӛO��\����8�{F�K��?���yTʿ�N�K-l��]L�p}!/�|�$�9�ϣڤ�]��w�Q�d&����������{r��֭��ǜ9k�~��)� S�b���,�(/�	��{�V�/�w���X|Ǫ�g+窎g$��Q�u���=O��<M��
m)�����;�1��k)�Ƈ��2��
������V"��MϨ�Vd�\�������J����%89�>�]�Yx��^ݮ�j��U�8��F�,���[�.Yq~9���K��t)�b�zQ���ׂ5'��'���]�UwkVK��+�$��q��V7=�rA~JB�
X@�E>�?�Uojĳ�P�:'�W��b!�'�g���Mx3U��:�����v�*]�����?�A�xG/��S��b���W�7~�EL(��.y2�ٮ"ؗ���Ƒ�ƩJ���+-ؙץ��B�g�z� �:�� ���X�����Sҥ��6/��x��W}�%����u?�<av2.�h`�M�&�d���G�������i�T�\�I~B ��^(�p������/�B�T�H�r-����C瘈�Lr�(E�R��{���Qc"�� �n���|ݬM�ȕ�`[�2��2>�KЩ�I|�R $���mqvN�����Jĕ&��6VY����a�f��}g)�7h/���%�(�
}��=>��%�V����/T���;������]訢�O7��*T!���W\�-�R��I՜Md�33y���Ȍk`���|'��q��케}(یu�������O.�|�~������`°���1p���6��׸������>�F ��=I.V�2�M�}&����O0�������8rY}b֛���#���h��/bi�����jc�0�XBE�14� /��Q���4ډ,�����E���S�3I.nr�F�T���>=�PL�7�#EvU�к���єt�P����up�yb��׸�{ʰ�鏺rƚ�k �kxZ���o� �k������m��a�)����J���)s	gq�E�����1��DV�vxp'�qƦ�,�ouk�۳�76a��G�Iۻ
��O�;�E҅�-���+�b��K��ps�󃬞�+�,�2,Au�
a��S]!#�S��` U��%�f$�u��~P��N�[� s��'����,5���´�Z�H�N;�ӔK��-����g�<O*dob���6���14a���K�����&vˍ�!l1�C.��Eyi�N��>p?��(�C��1"��P���ȭ�[O7z�G�@�]h-h�YX����M_g@2�ob���c�.���Xk�8�����#tT;,�>J-��c�a�.��q�D>A�҅zU��X��*� F�49ר�^TؔI���5����ն�~�z��<�����C����~��+l<T`2�|�F����*��&b�f̰d]`]`v!ZJ;�R��L���#�l�G�������������]o��)T�U2��N��B�U�-�F��~��������w��c�rU���,�ӊ �1�g�f��I/_�A,�&��JfML�,e�*[�5AѶ���dJ
~���H�06��>Ȱ��i�6��1]:�G�ǧ���8�Kg�`��A�=��/�q:]y-pP�'�i�E��>g��NM(x�I��)I<��!�<,�J��w�(v�b�s���f."H)�,Ru�Wu�~~��ܐ�����p�h�=_��6�������m��B���MN�����t|����+����$Ld�=���/�����)��yX�O�Gޗ��%�;�4m@�ZM�'h���=�7Q���M�%����F.�E���b��+1\p6�S�2Jk�v]앹i��NsB��7�s.�Unţz��Ck��E���jW0�[ c2�4�n)�g��6H����|{�ֳ?U}�(0���`����;��ߚ#^�J'E-�O9%~����^�2C����ѱ�f?tL��r����W>�U+^x�[��kdk4�����c6��=�䬅>���:J���ҳ� �0�t��fd��l�Ѳ����"���:�MW�6t�	��������l�"W�׈ r,l=,$��ߪ��і�����GY��lnp�yx��W�j�=��zf�O����K9(�9���{��ԭ&�Ũ�,\����$���EM>#���y��:��bml���L};����/�ǥ7���)�H��3��K�JM#�����<MY�D�a��d5�����XfH�8�C����2�1��t���^L���WNȾGX��I��Z^_akj��������siKn0�D�[g�j�)�W�8e��!h��|�⁏AE�L�U�'nK{��^�ܕ��E�+qVJ	� ����Q=������@�UO���xE)��^P�6X��j�y�ۚ�����s\�i"��lI���9s܊�P+|y�Cs�j�ԯNC�0�g�&ݓ�E �xm:n��A��E��+����`~�y2x�>~��{7�������D�DZ��[ú�|nH,����B�
�@� '����۟�7�AX��e6��u�dIa�Th��^~�ج(MR��Ty�n؃�Ԅr;Ļd�	�~EA��V�A� (DÜ,G�˹���>Qr�ej��A+�~J�Us*���"mto�9��ޣ���(�ۚ�c}ߕ�~z ���_��& hR�4����7�����>�k�)���,�cX;n)��]F�m�`r��6���B�@�q�_�Qk9�*� Ww2��K����e�1
�96F'��Eim^E'�B䛒�b��bE��N���Fd~�>] m���ֺ��\P�#���/+�o5�2TS'�z�Fteb����1�PB����M��a⸤N�|�bS�`�r"��,���S�u��Y�|=3#�',�=�w˶6��<0Ez1�W8��<E��J��1�]�?v�\����d���z ���.��0��m��8�/��b�%�]W�R����^������ē~�UE.�WT#@E��/K!�>bUY�دQI��=�=�N�VAF��{�h8IĹ��U�w-m�����m����	Pލ8�2��ݿG�Q���
�q�_x�u�z*��wF_��]�n0�EW��U2�s�2����<��TI��жƆ��w�y�Wk�j�p{���a!u�C�3O]l��N̘��}�-����0n�Z�t� �ythr��e[Rv����b���J�/��P�FD�ސ7c���E����!ߡ� ���N�4,!�Z�gO~H��F}�ߥ�`�o�e��b.�
kY/�Y��rw#�y���f�V	��92�����4"���W��ƕ"�'q#3{౔enT�������ws���yY����a;.;���1==v!����哟��$��puf��
^Jz����y'�}��m]�e��dn�R�*����KY�S�a�=!���;���dOAb�?����\T�#�.�X|�"��֍$ֻ�13e�D��,�Y�YVR ��2�c���=ފ�æ�T�YWv�퇸"'��6�Q��yB�kF��7fӥ}��P����>�ad:W������p���G3�S�p�@�]���-.̑e�`I�5s$�g*�b%�>�z��6+��@@�3Vu��W�BYU� ���z��g�Y�Ч�Yu)�"��Q] 8��5wY<��qt �=��KטD�^�^k�9�IW,�[V�������|sσ����{�ݴ6Bd!3�I��Ev.�OM�{g�Ie������+A�	C�����
�z��v��U���g��^��1�hE8�>s/��;���~���s��*�ߘ�x����}�з�Vs;�I�OYx��MJ3e�ep��*����=�W:Ȕ��G�.xm��d��N��r�7d������[aon��~��H��a���;�>p���X�ާ���Eo�0%/��w���_I�{i��V�%js0P~��2v�:}�
��A4�10Mb|9n������f��9eRK���v	k�ť���n��Vu�Z��z$u�+D�ֿ�:��FK��cV�K'�o�h'Ԅ*���b=쳴m��> � �M���?a�m��9b@�ŭL��q�[�Q �/�I��XN�;_�(c��]�[V��W]H]r�]�Z4����:{篽5�T��FKGduǞgE�q�!껵���6G�fp�Pb"��ɮ�tࣲt�հ�������%�KT�QF��V1#��;%��k�!�ľ��~z���6em*~�����p����ox��&=Ძ���jߪ<~AUT�j^��{ư��)�1j�Lv[�S#�>T�Y&��K�Ө�~�|�j.mb��z~�f��em�u�x
KD��ܹ�M%�c�y-B�X7������1ALP�.����2����������覎��6de�?F�Pe+��*��3��\��������i_��F&�[�N��1
���U9�y'��7:�\ոW�Ax��
�.q������ق���؝�A�����g�l)+�v�aF�@�\A�5�D�t �.�i��M��;�t�uͭ��kkϤ]�>4%o+d$|U���˕GJC����:/�-����_5���C>R����⦳\�I�n��G�;'"��D��F�5Zk��!��?R�tXqBn����ӿ��Ǣ�=�(� )�����;d��x��|�S�,,��93��	�%˦��4_��v?��������S�s�F����J�\��j9��n�=m��d0�e� �K�6��'3��ϑh�*��r��n�z�oB-�:�a�%!�v�c��61�&ו���Ȁ��˂ޡ;����Wc+'Kd��}�c3� D��"�j��ܵn���H����/#�?Cs�/�q�Ys�g&�N�A��`��E��g�r�o��������?K,K�m�7�	X����;O�C�'� *=�S��d���%+�17�������5����R�D��H���Q>@���x��H�W~xذZM?R��86Fhm5�sB�3)�%`�W�Մ^����C���0T����h|Y�pw䑜Vj�,IQ$ w}���T9<CZUxz��ԟi�c�w��~�.�"�$�^/aohhd�0�#�|�?�&ȂqB�-Ů`�=�z��3}�9�]τΜ�MOP?�T�oќ�)�'dk3>�?��4�U�^�#
up��m��� Wڅ���T(�N��8���UN��V{��j��O&m�O{����ʇw�������r��F��W�>�B�(1�l���� ����2�	�._�T{;�9��u��"Ď,B7g���O<��/&�c���)����;G��#FS��͠�[T����#������ڑ�E�3B��B�B�,;WZm��������.��楈.S��ŅP�@��7S'�`+0]n��O�T�%�W�Q��6z
0G��{���q죹Y������u�A��Z�Gj)I��mg�=��qA0��P�Q��. �vI��oϵթY]�����>NfT�ٿ9�m�my���3~-fя�
���_�?��l�N0�E�<�	Et�o���b.<�M�m'!����XDn5��l(��C� �P:�_���f������?J$$Di��A�Y���3����	�=��[i���#9�X��G�����% �w�,/VW��~	�������V������7���Dd�'p�#��i�L�m^2:gW=��-���2��n03�TY	��G�n�g,�i�`�W2�:����`�H�簄���tE˦]�b������u��yς�C pfҡ�[���\��7H^)ќ��]�U���7�z~��Dv*I��y��Oq�����Mm;�n?��}&2���i�Æ�����k]������Yi=E�e�$քT!�B������b{X�>�\�0��_F��u�g�jI������LRQY�%Fx�������k�c��wF9�&�M��`�f�8-snr���`u �����d	ݐ;�Pl�	5�\5�5'�ث����"_΂niO-������@z_%���_�b��<����?�I}��~{�"��Q��8f���'`�·�:g������Ci��]A�XV\�]�	�i��_i��-�����{	$�g����9����b�0�����X�V�h�C�7�㖋�Q�`��u�Y��fڢ��ol�o$����_�<���2���s�x�t�D]�z����Ţ�{�=�W�P��]�,JW��yb�2��/�9NX�C�a��FS{����Z}n��fOU��6��z�@����2��kLe��ۨ����G�N��@UUyJ����$5W���6�_[ZF���y�p���D[��U�+I
�y��=���u^HԘB��H��gt�S��e�:J���U|.U������	Cdl�����#����x䯷q֎�,K(*l�x���M� ��)��5�5�=�]��֜����<�sE�o��*��N���1AN5��#D7���f�c^�r[����4Х��m�~���Jٛ������#��0�kc��x�lhGs�Q��wɜJ�f�%(�*�铡tq]Ǎp���D�H�͍ ���X����/�p�����g��{�i� n0�[36J߫�S����4� pK0�w�jw�̍�,�0�<�(��j����E���W#�?���U1du"�J�,b��+
���r8��P�_�������_{pl�q!o݉�^M�_��r0N��p�X�A� ι��,�T����s�?ԟ"S0V������,K�\p���(V	
-�}���7�N�(O��,�<��G���r��f��-}�IHy\62 �%��I����|@5rȞ�6��ˤ\��V@+DoI#�@������V��!c]�]����(��B�� ���o��e֚�y����ll�A(H��"�m'��o x���ҥ�P�H����=�zT�Rsg���r�~��i˯���<:s=�P��]�����i_չ��	�ĭNeE(��D��t��R�59&�'�
���7�j��L�)H��s�FB���Z�����SM��� �.��ê�{Qu�%�4�a���Z�mP�D����&�� �hn�Ƀ��U���h3�ۇ�e����(t���[p_��x�=)ڿ!'5d���CȣdQA.���������n��(��DI*���(����ɳ�*}�Z��6;�(eľ�h%W��T�	�΂\/ �UM1# ��5�˒�%Y;��qs�Ӄ!<��`�p~����~��{4���]����O�B��s=3��*?�ѭ	��?~e�����=FьBf�o��M�)���ޞǐ��˄���p���� rO-��_D����r�wmZ�}$���q���ם&��_��p�h�<ʳ�u���bx1X���/������a>�@ϨZ~������n5�e5�	ȩ0Յ1c�q)w6g�?���q�.�3�,Q�52x-z�w�ԇ�j������ �y�t���W�-��N��܏X��֣߲zj@׷��cNj��Fk(8��Ƅ�0�!F�lEV����T�3�^'x8轩�?-T�Ȑ��T\Z���Th<�{x�s���No����k��F?��|�D�B_5B���2\R���{i�C����x.�nፌ�=�`�j'a,iu��`,�򱁫��3�f�R����\ݓ`sI�!=�O�H�� �`ڊ
�B���g[!�v�#���	
�J���k��).�i1騖�UCo��O�z���H̓��+V�`ɝ֥��q�}������s1(I���W��qR ���p2�4�o���s��X9e���X$}׃;@����&��f3R�l��	�����I��E�W�{g�si+V�g���IEģJe�!V�߼K w�D��к�I�9Yr&���Z���X����0ot��1U�/d��Z�JC'���vg���7!�{4h1��z���giTz���*������f� �ܾ	=U�b3��ַ���b$)>�۴V���VR��_E<�D�]�
��:j�X�C#d~ʬ�:���*K�~��ƨe���������_,�CMs�*By�=����3T�9��`����3u=�À�l7t ���S���z��i��e��"y�=�._5v��#k�'�����_J��2�&�c@��]5���j�W<�������e�6vI�N��ij�?am��/5�ACJL�K�����q����d�l����X �l�r��]��B.�q��m�<��i����������*�wVF��0����eb���j��Pr<�3�M��S
%� ��P�!������z󄍠r�<�:d�ç)p>F�=�pV����c`�G�4G�y'3����LU!��/ONiq�Ů��(7Լ�/2���Zp�ڛ��gc���(/�ҙ��A������|#T�5�7��fbd�����L �|�������'��%h|�]�~��E�����l;�����P��vR�K���KiS�%�21:��1Q��7�B��D���+�ѧ&��EGjt����� �'��=���Zݾ�'؟�!��m��@���qGmQ�
�y�{������gQ33*�nep%��I�[����C�L�'g��Z�~�9�)��$u?�(�c��V��MXJ:;pd����p��='���aJ��.��q�m��We�i*�$i߲�n]��IbۍW�G���u`�d�v�0�� ���=���6N`θ�mJ���W:Y��]x��q�x�I�*�h�P�M,b=]9�����"֣����y�Ѓ��%p�K�D�����QGi��s�7ţ�]ɦ2�p���cA�H��$��7��q!���>gZc�j���u�8���P�|b�u����n>��0փ��p�2=t4>���(d�9.]#�p�ٸ؄��S�z���+�-�=�N�Cҧ�>��|���Ĉ�4��� n�㈕����He�{C��RzP&KK���J}pm��&Ҙ�G��RF�\Q�Y#M�E�����4o�-k2q�96Fb��'S�J�꥓��Q����.c�%�����Z6����<f��V?%��zUi]4�ᯫ|�s����ғR]�Q�?��K�ѻ�G��?n���c��]e6]L�*M:C�K��كz�}wCa��[�ғm~u^}�hY<7�bW=����F'E4�� �I��K9����u�+D��9�pyQ6�͡^R^o�G>��'�'-��58�س��k�26;w7`Y��VvZ�����z6,�,��
4�FW[�b����y��&�\�Hy9�rv�߱�����z -PGt��	<_�G�s�*��6�gQ�5����Tqr��!FY��@��/\��<�k��&g�/��-��1��ͦ��o٨�Y�!��T������t]�I]>���З��c�X�B�!x��)�{��9/<qv��� ��}��m������'�dO�|�#�ԛ(�"�;go�+�:C�u��W�����<k��wH�楅"�r��ʅ�Um
9(����h�s�h1H�SŞ�b�E�/-���R��EY���[�I��D�T��71�@mX(xf�������}��jOŧ�8<rG`m�����߾1̼P����Fl$�áɐ�,����%�A�=*@M�Gï�Af�H�GYV�Y��wE ���|Yk:ԘJK�)�і_#���*FS��_���E��[o/�w��{� �lPT`��X�P����n�e����5C�(��7�JOӽy�5�㤮$c�1����3�6qn�y�C��t�D�d��lp��SXA�'�$=�V|�d^4�'�
��/����ltB�^�/��z�N��+ad.�v������5���e����˃a�Dq�~�2�l(n^��z7��wyk�F� ;J�	"_���~����-��Ԕ��Ey�@�s�>�;VX\}U%֘�ݼ�G��yoۇ3s��ci=*�>���~���$1��;npW��[�m+�[����<��H���~nvm?�	��>ukL��V��)+v��
���׹`va����Ik�޵^��1�"�����fl��A���_��xR�T\,|�a.!����V.�>:E��zm��t(�9��Қ�e˹�@�U���11���Ə�������*1���:�50�^�L�=�v�E�St����Íc�5Zm��9�����L����0�q$ɕ�X�}�_�9��D�֏�W❣��'��^�0���1J� B�j����[Z���.�cYC�>d��]5<�i��C�_��-� �V��U��ߗD�?E��Ъ�/���v�|�G0�����9�ۢ=��K�3�$d�	�÷�;]ٟ��k�1�q��.o%>�%�d[[b��Lh2��G�V��N;|��ݥ%���%�T�{E�(s����yb9�:�a�OƮ�����o}�XD�V��V�v�g)A�F�ݮ|�=��~d�c<���P�X� ��_y�_~���xv�")]!��oxǞ�d��3'���z�l��m���<)79�V�]R ���� 0��7��8ş+�E�#{��U��9w��5��+Rҙ{{Cݺ%;�V��`�Pf�����j{�}h(��r�+l\G|&�r�w#ȓnjݩ+pm��X�F�l�c2���1�*&�S�h^GW.�^.̈���:���]e��Q��	P�P	�����ƈ���p���#P!s�x�� ��:��[�fs�~���Ȋs���'(�L���_�W���8驀���#�"�q�Nc.�epɱ�"b�^J�#L�Ц|9@�$6�Y�n���L寧tZw�`N}�}�?r�;~J�ɜ��4���
EfA![��	��H#�67��8�A�b׺��?OJ�[zi������aO�<GM���v��N}�S� _Q)i�\B�����d�0|�EEU��"�Z���CC6���*�ܺ�r�ǳW�&��a���6:H��xwt#�9�b�~_`�J0���Ga=��B�r[ ݒ�@9|%��d��S)�{�cR�JYW��nG/Ė�Y�~.e�|�w�=�+I{|�}�̍ {�5���PP�	6U	ޝ�F͞i�uj����ރ� ����Z���Cf��b�a�w�B_=z�Y�a}+�� [�X���Ec3*Pn��)�E���6���,c�$���I�MW���>i����9�n�40����|�;Ԕ��V�Җ�5�iq�6[���r?��>���]o�����vC�+ų&���D
G���ߑ��j�}y�*�ُmn��>t �@�5C��s�7��O�?�x�m������s �J�O�3�&ږ�e�Ț�'S�����D�sPW[䳣l:0��Fkq��\ �S�<�WhH�J7M�a�2���m<�l���x)]%�t@7��L`��$ƭlt1EO���5�}�IS�8�	D+?oQ���Ƙ�2pg��pr��%I��M�uªK����g���q����m��*��Y��T���O���^�?b�֋f6�$@~x��Æ�n�Ixgj!0Q q]L�)�
]�&��/�_|n�_���K�D�i�_�,j�l.���m�]D���s�/_��#Cv�ѰF����|�_�\A�01o9;e6�vG�ѣsҝ�(V��D ���.����]�������$����L#���^i9V4D>�y���L#Έ�Ů��^����%���K'Y�p����`|��0*,e⇆�]KSP�,|,�����Q��X�.�'O�5��W�c�c?�����;Ps�w񡁶HI�HX6����d��w��H�Ȝ�m�T���؛{h����X�Ťč�#��e����g�3B7i��J���)�ǳĦ�ja��
�̉Z'����A��*{�M�����ʻF���� �Af���ж�N�2�r�o'��0�����'��	�e()F�K��#[��4�K���B)c�~�F��&&Hs^g���]}7:A$���w
Dλ$�+5���H�������KߟI�I��f�u)sV����&1�X�
X�]����%M�
|*�i��	�mj�x�3	��N`(�ZfH�)�gq��_įf�0�����:���d����{��r[{X�	W���*�a_���ݣϣF�`&����c�H�(��{Ju�H|�Ј����t��@��h�m�t�ތ�_b�[��Z�%��`P��Z��/�7�M�.0�[�w�C�q�D�ؚ��ng��w��Ӽ�.�7c�-��T����T6�y3�˜$	وʝ^�"�	h�ns��:A�'1���(�_+֧蹩����ÇѺ3�-���'�|�o�n#o�+풞2�U3��=Q�1��^��H��ƮV�k�A݇&��D�U��7�Bps}��:�c+�O�(g��o�۔O�������7�@r>���!��'�l�U�(���IR�ov���I�S�{����ҫIE��7d,=},�˿;�:���������> c�Ϸ�=��8��ģ]Z���l�����9i�p���Mi��C���ƛU����چ�,�Z�A�E�.4��l��F�Ȧ^��$v��
me�_�34_mE%q%�ȴ�b�P�x�o!Ar�S�m�aE$�d���RS��H�bs"e�6��>a�����o�0L WJ,Mh"�2|��;*g��2_+�<B5��ɫYx0�VN��ߵP]aSW퓥5��J6?9��+���P�}D�ؚw�yj�<q�`��	����KՏ���&Sz�D�<'�L��UE���/����%�R�T�&mU�}�e�������*p�eC���|���cu�ꓯ�5N��ߏ���]WU۟�����P���g�����a�����8 �l	/�w��9�8~l�"2��{&�q©����}Ϗ��ޤ\ZM	ܨ����Ѧ�� ��ӧH��
��G�� �=r>!�~����~�@1;e������(� :��
�F>�-�h{��Ƕ�qT\fή����	�<��o����'>�|6<at��N"��N��bk�,�=O�$2�rd�2��{���<�1���>�#p���1f��ǎJ2� "�х���$����\��C7	���1Z��ұ#�tԗ�&�L޾�6X�"����A��+�@��EH5�1D�����(��s�񨰐'�ۖ.�s"]Wǜ#SAIT�r����]�9�v拾����˺\,t_��͡|���Ӄ_�[��K�t���E��
�	R�Ǧ���xzŷ���5���Z)8f����c��i���~x0�T�-v���l9��Px�qQM/N8Q��k'�̔�Of7%D��t(������:,A�ٰ�?9�Oz'ߛ�3i �>= �0���Ec�Ө��	,o���z �ʚ��ˊ��N�U�q��=�bx������T�R��B�=�J���y���亂����><c�d*�g`�����}۵��~��H������D��Q�>F��]��)��K�$ũ�U=SH�&� �}��w�chԣ�����>�d�Y��r��$3�f�+oݶ�+���h��<�h�!��X�9푐Q,�����o�f��;�V|��0���K{�����m��`�m��U�]�>�@�:c$�nF+E�����h3 8�|�u	�;��vD.�(� 6�������X�&�pfb���c���쬌$_,B��xI"�N=�V?϶2ߋ�~(���W΅���p�oHS��[�B��$3�},@�����d�ce��A)��r!���7 ~<���Z�mWcg#fč�k���:��8���I2�~����km PX�h���A]��Cj��Y��������Q����K§?��=�M���5�ߌ�NM*m�<v�
^z��q3�8x�wc|�5��^B5�1đ	�LKu�rBm[vBbS�.��3��j���:�\�q^$J�X�:	�I�r��^V�p��{�Z�l���c~[5`��K^U.W���RO��J�6���a�+�IE"���@	`��@)K� ��.��TH����5�0,z�d��L�L$�ؾ���]43�᜸ǜAb��`�,����&�����N�%'@=��5�Vj�����������.�k��3"#���Φ�0>5b�H��c�AU�9�y�ƴ<W�������mJ\U�N�l=�/1�z���vv��8��&�]�A)'VZk��z�p�,�/ ~��C��Y d��LT&f�;@��ϛ��� ~��S5'��p4O~Z9f�皢�w��:AL��E���d�/���lf`˛�,�Q�e2�(S���o������_]���1P�hW�?kNwo�mb�jb��&/�戂��
Ɲ�:R�V�	�)�,�R"+�����m�� ��@�	P}��0���IT	�iӀ�KϴĤBa��-����Ҽ7T�Ox|��~!���
s@c�FI\��?��'�ϬY�>��RWd����nok_���E�zz��~eZ�����v4����cD���=��h����1��5T`��H����(��c�)4��'*���1�@c0�#F ���prRY48����\o���.SHl�i��Q��$���DcS�N�����{��j!f�r����@�P"��N��뷠�;$u���G�rcjR>��)Q9�5G ��4��c1;��n�?���	����j�>ǥ�l0Q��_̵b��Oh1����/�H��Z[��Yj�Q�r�⿸&�䧹`�\A�-����?��UhP�g4_5ӥ��X��soRA�Z@5ڲU5��J����6�4�ϐ!�#�j}�=tt��� �����9��,���Mz
V�������HyD�cx�d�+H��y�W��7m*0���>�<9�݃���<J�]��lߞc11gFr.]�6X9j���Ú�G�����c���	����\WJ��Rb�
z�#��U5s'�ڨ�r��!��.��l�_�V��q�w�ր�N� �i�BdW���� w
�*Q4��2������Q�w��D?�f*�>���R|H�|A��cN(�f�E�8��PO����-WSaԏ�JxvM8�F��A�/���Y��v�����1�	��W�d���v�8l��T�z���L-�����E�Z;苰`Z��I )�̧�����J:�pQ�ZҨ.]Q*#�B0r�_yǪ8d�L~F{H<�%6�[u{:@[:��� �lSC�|$�dbh��(��ͯ�]��S‐z.Q�;���9Y�,ŀL���+�Q��2��ԭ;V���1����<_�#�l>���|MW3��Z�����o����/��"P��һ�u�6<zw#�e�9��Z*��ڳ�#C<������)~X�W��v�L�`	QJ�֎�j��*g�w"����r��t���%E��C%&y����& WJ���\
�����T wt[��z�o�!O�\,��r��Ty�{�z�ۀ�O�V�I1^ZQ��N��hi�B�Ѕ���Q�Rv�ڌ����0���棆�P6<�f��y\�'�'8�?5rP��:wp�"Aw���٬���TyX��<�{o�U.#�iߟ@J[�X�!�pE��؛��_�J.��,�hx�/�+	l�����=����
��T~^���p/6F�p`����Ü��#Z��Ӑ|��9$�.֔gS�s�U�c��Gľi�d5?Em��B
�i�F���,d:� ����G+�i��l䘴gMgʅ��`m�������&C��ór<�R��M4�^:�H�x��1K�n�M,8�������翡|����n*;��#DiQ՝q��{۹yb��֨�E�nI�!8L ®�Ⱥ�e������YR1�G�W��a�VRM�FI�?��t:|5=
����8u
����n��W���?t���=Yv�W�u���y9A�V@t�S�k��ifk%_%��d*;�!H��3��`�E~��״�w�{ǺR"ذ�{q�YB���s��C��a�6�z��y4���S:�����-�|W�\�L�뗘�P�ֆ'%;�A(]᱇�J0:�r#�+��U�gt�������Id�`���I�p����A��@��Z�}2Q��Q�)�������[����G�p�9�LD�J\+���hO��OI���Ί1·*�,�f�X���cY�}�߯�j���<pǶ�`+����|a�;�2p�:$��L(8wpN�+c���C�t�MSt�����Bj�Q�T��J:ط5KI9�6gĐ D�8�؛i��M�N@��|	��Ż��u�-&x�+0An�%��l6�e�*�؏)C#56�EK>T�u���d�>S`!h�∟5/:�}�僐��v��Y}
�6�_Y�W���0��=ѕj�)�A��*sY�ze�6��	6wި���s4�܆\�]n	���R�# �f�ӻ�)��s@�<�n'�bx__��7+�����u�?`��0ae�h��䖒��0#M�F�Sw3�/�����ֹ��GCq�w����W��S>Y�5^s��BG���-��5ؽݛ�_��f6��#=�g��C��X��*���=�H@�w|�9y�Ң���M�~����=i)@Q��̫������إT(�-Y�ˆE鋾�8չn� G�cl������ u�P��C�� �|��w7���w��"���0WE��&%�����eB-�֕ŝ�����;� �f���o��+#�W������3��@_�&���i����� ����vY�A49���^��f	*��K�:��L��
O�9�N毥'��oئ��>�A�xp�p�u��ڌ��<�����c�B�5-|�|!z±���� �74�[z-��%������<>uURF
�'��<��$��~�q�8���L&�v$�ۓ�����k���?eK��bM��\�w����~U�3��cW1��yN���{'��Ƥ����He{r���Eg��K����6M��� ��JHY$%R=�Xj����{���4��ne��; �ɨ	U1��k) �LQT�x�u�ꂔ��}���nϓ�<�R-Q/X9 b��o\}2=k��Fl[�J�sP�nqZnS�@𡠖Kg��C�Xv�N�9tlz���q�e彿�<�_�/v@���r;4����Nf��;�pMƈ�X����q��lj��b���X� ����}��}�z'aBm#��T���IRܿ�t,�zo_T�	����ͿrVE����ϖ��]GA�����9��ٹ���3��}.#�m�@��4i�6|�u�xj�mGi�DF�H����I��g����Q[ ~�68I0�ag��(�m oW>�X�7�BAɵfd��E)Ӗ��	��X�q����k�jmh�Jk+�M�\(�^}ޖy�&�F�]Q��	��A#3���k�2TP��Y��$����P�jQ��b�x5ϧ�W1l%Le->�s�=l�����s���_����v��D�|r.)?����K�
�� ӂ�Z�%�}ًW�s4�	�0Q�������ޖܩ	n��K;ݒ

B��m(^�w��E#��p
˨ׁ�<,@Q�r�NK��_ 6���{�6�����@��ZUe?�|v?HbƠ1��i��Eˋ�j=ԕk��q.�c���nS�����|�H�m`i q>[ɠ��]HNvO١]+��SG�oO�r��'l9l�O��E!_Ѭ�`U&I<����Ȩڏ"��F?˵η?�j%���sk����H�w���6�]���I��J\��?�{�1"Ȯ�̠��ɔ��,��t&�|pPF�c�`	���HU8D�߰օ��.Z<B7��8k�k{�M�/��Jc,�]�r�~⿕��14 ���(yز3�v>#�� dtL���H͞_�9MŘ:�-ܳ��,'��$Cm����綉m\�;V�}�[��uʄ���w\����&�!�U����ʱ4�E�IIf�hO>�$ˡ�B�[�K{-�J�c�Wn+Rw{��kq@<}�@k-4 Ka�7T��ml�s?Q{h��;B�o�v��FC�_t[���Uag��D�xWz�+� �ꎀ����N�jh9Kg�휵g��DL+5�V��q���rh�@4?	E|2���J�RЛ��Ϻ]Ax�p�]C�����@j���E�cF\Q�Z�o��i����U,iD815ӊ|Z�/ݺ��ǟEn�G>��dfH����W�aAm������S�*��+��W�B��Y�x���P�ҴQQ�cڔ?5�,�7���(���GH��>��B����I���R�&c
��b:)P�#>��Ef���fM&M(J�/<8}����/�1�y2p�����b� );V3����������,���5Yn�t���`��)DWU޶y��Iߺ��3�l�P�X���H�6G�"�@k��ZL]�a�����A<�����Β��i�
��tޣeu�d )�ɐ��zaO��NJ>���P�?]�Ř�>V�e� =�H��_.�ÌF�l`�q*�ɵ��i�}$���:+v���2�OhF�%M��_D X���¶��@�L���Ie� �E�Ƅ����n��{���$��*} ����HK�_T��ۤΘ���(J�o�MMM�z�f��)��p6�k��� ��{J��uD[!s�1Ų�R-��A����+Kd�ƪH͔�}b��Le=�j���s�xL]h�V����=n�����k?`e���ݢ��S:-o7�����7	d/_	��Qc"d6�ѓ�hU7����1���Ѽ�>�� ��< �������/؋��{�<<ցNI���#��Ѝ��ҹMF;n���m����_�XN9!x���#g�3�k��Z ��,g��A��w=��:�<{$�?�W���γ��1���&�̨�⩹�H�ЮˇO0p�=5b� � �r+����8���i�����/쪿>`qP�%r�e=�wE]y�0HZI��R�v���'�%��?{?%�d�ӕP��]ۂ�-�8�0��0��MA���Ս:��Nf�H h�@�@yܘ���0�~&/wpV��kb� %�ܘ �p��(���]���C�vK\c���k�w����K��	�kk��t�e�fg맾���b�:������i��I���A�B�|��M��0\�ȶK�����<�M��=�|J�31l/�4��.�5餶b��ʂ.��!	�^i��n��`��>��#��~rw�9"�vIł�����w6� ]�y���C>5���dj^��èSY6��>u�Eq�ϛ�}��H�)�/q�T���P$�=�
SX^v�B4��IϘ��(1#�2�2k&��\�,BΜ���>Q1y��6.4�O��1L����L^����]���3wΪ� b$V)��ʣ�n��e%�yaܖYS�����Z�������c{�%��$�4`�U�,��đ��@�ώ�ȵ���YNW��3,]���J�Pk�聅2}��M�́|!�-�-S��\����5�x�}lY�[.�u>(���3=�w���Q������-	k�DU����g*O5.OW�Cx(��Y�=�>�4���cT�
��Y���yڌY��>}2��T��`1c2+$Ӹ���z�&�q9�.��o^J��� �|�y�.0��x;b��sm&5�-���O ���a�G?H��6Z">�J��a*�yU��g/��f6R֗:_����ח<���h�o8���a�~�A�@�VE�\�} �`U�~k:�	�c�5��8��2�ъbAq�v&D���r��7^�72L��n�~��S|���p�_z��"�[;h]F����2������t!
B�K���ഥ������7�~ę=w�Zm-swk����k��*�����eGS ĻĨQJ�����c�v +�^?诬d�pm������[Kq)o�sWl�bu�$0o�6�P�~�5�������,<��lw�1�mA\�$?��JQ~{�:Rk^�ƍ�ia�s��4U_G��]DG���`X�x��~�@��#CV�/*d
�M1,��:�h��@�)�-�E����l�G��q��-���RGa�ftuVjr�Om-����r�P�d������KI�c����M��#N���aE���.!�#�.�
@�kmt��)��M׶�����ʔ���\^��^�d�Ŧ˯�#b��]���"�(rsX�Y��>g�(煱gB�r��?�U ~T�~����F1��Fug c)"�Hp��m�~t�mr��AQb8� _	)�iʴ�Є��-��8�KN�|�Y�?�/�8z��qX��m4v����Z�Ӑe엃N����Tw��E�u��p�d�CRg:�g����{���W!a���4F�0��W��h�U�*����*�g1�VEV�+Z�3,��� qE�l��9=���a����n&���n"LO������n&��S&F�/��/���(��%.�g�/þg�즓���2F�E�҂x���i�,Ѭ#�!π��2����WuJ٨��eX���W����Çl����X��<��U�N@����E��e�)@����
}��d[�4n��9�>�zxO�z��b���v�yiïɏ��]�i(�H��&8��3�=���2��vH=�AF�UE&�L��e�{�WXxh ���p #xH��?a��Yˢ�b�<&D���A#8�Wa<��/v�!Wu�8Q�v�pAN�/�}�|,6B��k@[�M,�4J�S��'Է��!3r�M[�5E&}C�u_t�n$� �/@L�N-�r�����^ ݡ���a3!9Z��E����C�)�ڪl�:A�f}��S��%�h�{A@4��i�.��DG�avX�s}��+��W�|^�|�;�I��l�t�t��m�+��J}6Z|��t����Pep��P���;P9�g��������d�-�=�M2�=�oNQK6WN�Ly|1z�s�N�ա����m�+����'0��9P>�qޕd��a��o���C��l���P/�	v�j��J�-6A��w�=��n�,%�5�P	A�������%�_�#��G��`�2r�u����P�P9�gX2B@'��� <�;1�{���5%0D�,�>v��x�0�q4�Џ�*�|xn�s^M�?��:[��c�(m�L���1���a1���N�d��q?/�7�5L��C��=�S�J���/嗘�a}�޴�#�Nڋ��˒�2�hC�>�o_�6����P1*y���$��ݫD�γ��j�{������o�r:���L��8���|�5�V���AbupaFN������e��s�G�M�̵M�����NfF��թ`�ɡŠ��*Xݿ��υ,HC�N��h��$0�f*z�#�S��?��8��y�������>6.0������m91/�<���#���4$u��lo���qU4�Dea"��N�AU��G� �lp���?*Hw�(�Z-U�j��Hڝ��;�RA;�c�>���cx����l>����u��c=���a�;��oA���������d�n���"#=)|���VW�#2�{����T�_�p����Ҕ!dU��3(�o/�-l��p당G^���:^%�K�P9NY�n�!���"�{�Y��(�=��]�{&hC�~�omO����X5:�չ�C�y%,��O�/�n�f��Z_�5����V����L��_���uf��&��!|��{�բw��#L]�ǟ�ֳ��c�[V�e��?��[
�j�W��r�ړYƛJD��f���؜�,kp����U��)Ү�RC��ӟ�f�2��$P��)�]�K�<�ڴa�t�8 �nr!d��S�����Qɩ�xPIc��:����3u8�j���`���ED ��V5�䍭5ӳ�=�hrAw���v�"�3�!�܃O����WmbZ��p��#��1�P^�#1�_�j���Q�����

���5�3@`��N�ù�i.w$%��`B�D�]!��5�;۲'vq��s�[�r����X�)3Q�s\q	���Z?|vK^� �g&Gڥ�xb8�~������ښ³qy6j�y���}�����(�-����tYݕ�B�̸��(��$.ze�2��7�Ee��n�+ߘ�X� a���8�Jq.�]�����g�ѭUy�u��i��"�'D�:��,��9��:b���!��˟e�U�k����*��%���` �i' ]S$�X���Jp�S�2yu�	S��� �	w�Ȣh���gC7��A#o��R*�ޠ�?��S�Di��"b�����EV���l�k6 ��7k�e%����m�˹����^��@t�|�[=cj�z��ϙ�����|��3��}I�e��eW��\�)�ʊi!���I����%�Lx5ku�t麧��^e��%���0����i$�hiGvJcƭ��ֹ�w�Ld��Qf��B�Jh �x�?>m"�9��5TVX�?g_��*!2b:i���~������M`�Y�JȬ��w)���8@��O��>�2}�٠{�jF�FL��b_��^��/�&�N�41+k�"��C�S��)W��1te�����Gx~�+MZQ���.^}�4VE�3<߳��Ұiq@\�M��%��'�(i�m���yA^i^Ga�XRD}�n{�Ļ�E�q�=~5;+���6�eI��H�'�+�"h7�0�^`]�V�|�]��r'�|XF��])x��s.�\,4����ߥ�,$e�v,�5c�g+�*�<�:[4:�2(��J��pj�sD�~�O[��v�1
)P�fɈ���C�_����a��~@́��+y����5��=�D�0� �m��+0V��v�<z`��4rg��{�:�T?���9��mVhӄ���0��)���}�2���_���kVD]����|�zAQ�*�ۚ��p ��ӛR���Y�Jx��6�@��(�O��8�Rq�'��������k�_�ũK��,B�y��R���[��0���%��l���$�L����_-��4��ԏ`��6jx���.a�!�Ӽ6%jGb�-�P�6�o����$�2ҝq�v�n�M��h9%�<a����L���)�@�ӧP:�K
�`>�m�K_(O�Pq<��7'�8��Q���]<}����{
�:[3)��/�m<yo����������sc�JP���۔=	:�)̭�~'	s\8�w3�$q����T�c�IC�w��s��K$�nIA*������/B�?O���{�۽p+3@+<�F�����	t��X+.�#�A+�5nb*���e�z��o��cN3� �Ņ�Z�'e����,�^q���r�/�\%bk�+��׮!���X��K�Ou�?�^��)� QZ� �U��vP�ɪ�k��k4�m!ހu��/Y�3?e��A���>�ٛ~<���5ɜVEҥ�+'������DM��fI���Y$G�Pg�l=��j���6F��K+V8��A����Хb'�P� �3a]�3P�;eI}���s5%PA�-A�PK�~��3�pB�GY2���J$���Ń�&���0�U�M{��\�nk���N���Ɍ��2s��TZ�A��2��A�աe� 1���;�u�p��D�N=�;��Dݚ�I��1l+���C���+��,)�7��ǡ�V��?ІB�hۀ$�-񵨆��u.Bq-��ܑ�g��_5�s[RyT,�F�Ӱ���~�T��I��ƾ�I]c����´̥Ϸ��S��(�Wi�L�x��7�цj�~m'9f]]V���RF���=�Y>���#�51Ð[LY�R��k�?F7�7�6�kY�D���9A��d��اL\��e�43�\�Ͼ�{\��@ߞ��M�<�Ю_i�w�
|���F�����:2���s6:�
��p�0N�NL�Q>�VЕ;��y�����]k5bk��O���j)+˿(G)�S�}q2'��u �->�ss�#��@և2�Q�������ݒ�i��)��2��.=�q4IݥtH-�z �c����}��B��꟱�HV�b��'�F�P��{�,zV�!��.m��s�uW�v�j�V��i���F�@�,���
0/�B�BL�M�������r�6�Ba��`��;�G)��'VkH�|� ���BG��a}'ܿ��-���fg�k/zC���1څz�#���i�.��3|��=�X�ǛVyS�:��@]%m#&�ũ"�j�/���ڇp��}̻ �8�d|;���k�=Ĝ�� ���Q�;^�6&��6,��x��)�T��;�ω��m� X19�p��.���Y�yl�p�=9��We7��q�@[o�>�n3m��t�O��$���A>���?{��`'𡵏�t���� ����l-��k��e6��q�+]���N�DϠM���Ѓ�����k�lbN��b������/q�?bOg������A�+Y/uP����,���i� ��E�?��4t�3\<-��I�EC:��qᭅ�}�>�2��(�ټ�O7k����*�}G��p��ݝ�������-N�#_��I^�Һ�@0�2,��$p�|�٬P[���݌Qñ�]�z���h?ɇA>�,,P���*-{���僈�MނJ{i1��et�*���rڽ��E߾�}�����gh��@H".`-����O�A����Z*.a=,FF�_lߥs�I{�������l�$���U?:$.z�|Z`�_�/vj�,�LD�����HtM^B{l:_�Ğ+a�^�
5"{�^�a���D���gc. w�\c�=:��}��t�G�S����z�z���c9T\X�9�K����W���+]����zV�a�D�ە��w��P�2&�aڋ�7�������ĳf��>L�h��Mp������C�p�kb�;-��oS�l2Z�7��.3r=����� }_b	�(����H
������-�}(/h��
��EC��l������R'碆	*KX	v�KQ�����*!55!��ʹR Yik�4^V�^?b3�t�*JJ4�@?���N�g��"lG4�L�2;i]�SZ�X֡)������LHc4`Uu1W��i���=�J.>����<����5�����5�\�<�5���(�`�+�_mJ�����n��������I'�&��J��/�1��R8�ySOk���Rd�O@:y�
���Vb��2��N��ӒT���t�����r
z ��*?6��/��5�Oj"�/�`>�{%�D��t@��X_=�v�""3'��nq��������ןty<�!#'h� `���9�� ���<1w���m���n���-�� ��#��M��W�����5er{� ض�O%��HG7$Ѻ��~DzŖ��ם���3�~�������`<���3w�����S>�̛ܼ������1� ��H���n��;��:�ˏ3g�%� ��ڽ(c��B��u�:���*Z��?S�ԣ(��Ҫ�G�of�T�p�+�,�!�����e%�/�	�ǅ�jg�:T�����]B\�>|���R�Aɴ�#ivS&��M
 �V.k!j�ڑ઼��I"̄�#�;���� C㼚�:�G��=W��#4��Gx�����A�C��G�.èO��5�T�Vv��ڄ-.�KBE���^{�_���y;���VV�J���_�nc�ƭ�P�?/��W}6綍�+��<�Pd�L��m��=n)�fy�q�8|}���Fѫ~��BHυ�/�'��ן�p-�D��,���_A�"������ D�C��r����[޼��6�D[�a�o�^�_�f��
^��pO>`5st��/\��u���0W����S�寫�?�QJ�������-��9 O�_���?
��k�$�"1i�U F!�Ѿ��ߪ���e_�X�d3���f��o�`�[�G%�oSnN����(P_:�Q�j��k���:0������i=��������?�9I�{��M�b";��)����@t��+�%j��Ζ9��3�=7<$�@��֖$^�걃��P[�U|9��5�*�Ђ�$,Aɨ��|�g��QO���u�>���Ư��=��6S� p��:�~߳?J�<u�ʩㄨ�����+$c��{�Q.�t,oW���NN[�d�&���:�gϚH �͇����N^�M��`�B�:����ltn]����9��R�hf`b���P0?�е:
�l�>J}����>QG���T�s�Ffa�Ua�0C��(��E� fD�L�Ї�6q�%����榁��"<��$/�h����ٜ�xp�Xe+Z��A��S<��(|��6-?�#���&�f�~�C>BL��c�N�����8>�SS�0co��9g��>e���r���H��n8��:�S�3d[�Rc�_�0<a�Ku'�t�����1��g!�U�&��W=r���V�&��7i��M�%g�.a	zG�L��!���A�q*���Y����k���X��ꐴͯ�$��9�th����E�62�f�Ӌ������x($�ew$^R��P��$�����ֿ\?���~�f}�R��iT`��A�Wv��q����m\z�u13.�=�V�Ќ1�y��$ٽ��l�@�g����;Č	��8��^4�(xM���s�õ��(������Z����-n%&O	T�/Ά� x�p �5�e�%��a�F�&J�x}���"֗?Uū�,���ϸ��7NG@�n�`K�q���'��Fvxܲ  �g$.}��t:��<u6��zD��@��e���4�z�M-#B��u�k�H����dMhnz�U��`34̕^C������+tn��7Y����}�����S�X!u��O2I�#�m�LC�a^����&z|�������-Z����4LKD�d�]�Ah�1��3�?�H���A�4��{E՟J��z��K�и|�/�\{vC_ Y�%]:��w�.�蚵R��o������o�H���T��ޗ�^	�70���4 O�<?���a�y�Y^�6B�ï� xN*+yh�فf�6�N�4�<߸���?�)r�.K��:c!�_�����Qʬ�����R��G����*��Zb�����:��K��Q���0�Z1x���8UX<|�X�y�ΑۊH��tW^bi�[ȴI��m��Ɔ�Y�6�bX�1q�.H��w���o\�-"�ّ�D@u��f���������6�
Hx�[B>�~�O��Ƚs����Pnd�ӛ�C�c(�ׁ)4�h 9���*��O'��I�>�ѩ�����/�2��-�{C���%�E�g��Z˷� �b9��xm����
��:>�ٵ	�������1-'�KT�����\p��b��3�5��n�����`�<Aq&���O��O`�a�x:�-��8���1�6D���Z�����ZG�_^v��=jX�5G$�S\k�=uc�K��
��Ѯ����[Y{�4���]�6�`�נ4�І7����L~����D����G�5*�?�r�	Sok�aj�uՔ��yӇ�S�1�$
�2%pf�/��ZuBfw"�[�1���@���]�<L'B�D0�i�ُ���i���f��3K �vU�/�<F�4��.��)J6�5�Ek��t%���w���E%=C�R�Z���A��X/{�5ug���k^1�/�^�X5���)�U�2�I�^8�\q|8�&8L�!����F�e@?�i}�_:J�4���^ű�g7���q���,��3�d�"�թ��Gσw��%W� ��`��ݟvg��w���� ,S+�����FP�@�/������cei�Oˆ�wf�f�|O����������]��sC��(<�#w(�I"����9�&�雇�+�����-k�,��S	z�Y��+SY�A:H��t���%�F���L{oJ�w�S�*�5����L��l��#�
d�u���.�����@0��CA���h�h����8=���K0��of�[�冨��g���$h�q�� b��K������۪�%��P�Q���3�Z+�_S�Fm��gū0���ᱞ�vU �����6�v3���:��Ȕ���k�J)��"U|���R�vK��r����&�Չ_���T9��y2��'����慰����]����&̪�S�W�Rx��������4lɄN�p���(A�H�r�7h�u6]�k蝟t�T�|�̭��k�M7K��������x�uC��/�����ݲR�9 H�DI^�kH��[�H.�"���Q�h�����+�Y�� �����D��e&ƖYop��}�6E��������	} �? ���,7I�����b�a���Y�,[g���^��������Yme���1~�GRO凳��pm��/�Z������K�9o�,�Ӭ�0t���u��Ϝ}v$�b�K`T�i6��?�ގ��뾜��� �xZD?O�r[�n��+��D�0[i?v�Cnt�~�_&��o��+��${���"�3���,�/�����ŵ��xq��(��/�5t�)}̻k�<�TWȦ=G)�eN�|nr���T ���٥[�F�~+{q\v��4��A�F��N��.��l�A��念&&+�v���L5�<g�i�2��Γ��O�{ABj�����ʔ��ϭ��1�P,�%�pxlFm�W����M��wz��t�=�d-//�t�w����W7;q$����v�meޥ�!DZ_G�::����N9����ߤ����71P��GE]���1؉w�5�����p󓒶]��:�J ���ϕ1�x�	`+8��2m��Μљp��d���)J�~M���)?(��p!`�]8P~�fz��3������A�^�i�#���Tt1���F�Buu���ñ�Z� �����$>�EX��0����e�`7CZ�c�4G촀��R�(��o}{Q��-Yfh�Nukn�$<0�//%�(T�_�[׬�=-��0�V�v(�m�԰��yY��&�y�����?��J"�y�B
mâ�����%̧	A!��nO��Hyx���͙�jP���fb�*�Ki�I+w��X����3�u�1E�?�|�P��
���;�;�0��=�m���ea�ne��t<�͢0{B�����w.���q�-WsT9���J�0�����ON�X����������xgTG1�0sxT�)��"cy{�\��s�М/[��׺V�{d��Q��m/;�J���kU��>$�uj~�Lv��q�|g�Qu,T��3�%��d��N	��U{H&�Vx��a�_2��>�J8v@dk�Fg�k��l�����p�I�=Ha./t��^�x۪����g��@��T�^UUlP����F�G�h4��u8��E%��ʃ]���w���qF
��7��hkNQd�0�Hr�,4Bg��"C�_���=��&�-L#��:�r�����y���C���UpM���1��4��<p_��������e�gLG��ȉe}8��P�}�Kܖ�Z��T7�ۙ�bm!�]�m:��Va`]S¬�[��$o�͌�� �}������� �.@��\�<}�C��0<"�s�˖⮬���E�/ZabZ�\Vy.�$ck5�n�k���f{U���,�mt�}�y��'=�ͩk\T}#P�`�QPr�"�[(���4۠lJ;x��3�~wS����+����W2�+X	gY�6,q����ȚC3����v@Y�>���6�S'��
�qG芷fu�Q�L�I�6�
-!d `��ޤ��vԝG��c�8ӝ�sW�Kĵ� w�� Y�v��ehS�g(	+��ﬗ�J>vn�
��M
ǅ�6D6��/��R�h/�L�,���|���W�N^w�2�0��Q3p�
��L<A��x�KH�)j16+͍�����0�*�um�6-�D�)���ts��n�t��[B��ƃ�@F�ӭ|lo,�yv沝��DD�ﭑ�[�jDƔ�:``��r���IaW�O�D���v8�^U_.~�����f� &"S�X�5Q<�`��U9�1���>h�����6g������-�������;�X��]�@����Y��}$�|,~E����5�������屘k�@"�6�R�"�PΤ>Lۤ� ⴃv��ّ��Tֽ�����P-э��X�⇘Wk~2�c+�b��!#�xrq�����4�!��66���Ll�v=� P<w��D(l��x/�g�!��uyn��0�g=�]b�������2��������ϭ�э�t}zM�T��L�2��Z]ԁ&�sUN����0Y��B��.bY�w��`�p���D3���!(2�%a�����{m��'�θ���!�/��sP���� :��A{�Z��kk؍��J*_P:D��P]�)�-%����9�~�,uPнS2��K��������l��Z��#��&��x�t}=��ۧP�~�F�6����gHSgϙ�*���U�R�L#�o:����!1���Y�r��k��0m4=F��DZVB�<���qO�tb;:�3N,���}�D���A�%�������￱1Tv��mQ�D�(�� ; G(y
KH2<�Sx��l5V�+�h�m�\�I��d4���r_�J<܁[�Pa-c�#�Ĩb#�t�]�)`��.FM=�YI�dj�XI}��o�Q:n5L���s�Յ-�/'��"{u^ZP���_���kC�+
�>�J�X���&k��F�C[�5�̳D8��W����^�]��-�u?���pU���n�E��T)�&*�:>w9P�W ��\Թy�Yh�>�>O
���� �n�mwMrv���#��r��`UdfKO�Ǉ����D:ӷ �2M��22ѵv_Q��Ce~��s��D΀��ל��Ue;~���	x��E��NŹ�Ju��� z���ԝȔ�ވ[�2����dJ�m�{�QN'J���@��{���3�9���1�U���ele�lX�rs�S 2�U����?��N�) ��J���Vֺ��`�M��K���D6���b$l;P#��:�	���6���;>f���MY6�5�ݫ^UP7��N�k�!fC��
?���{�m8d�]�a��*#�|�
lǒF�ں�`�YJ�QL(�+�Xk��C������(�-@#��1||����r �=��$h���xbI
K��wE�n#�Ө�S�rc�XU�]4�O��E�L�$0�`]�g\�;�S�{�kڙ���#�-��`����k�H&��"9�J�>kV���(�o�E��OH�t���K�\�?�0E���
\AĀ�7ѿ��@O�ӛ�VA�r|=qꓞ+қ�����KAbrє�HH�|�S1�J"+�h� <X�={���� �"�2�
,���h)�p���ē��;�b� i��le��s0F	J:
�#�T����-�w��^
�	�{��̚]�_�������p�,tp��"�E���|���|�I�AY'�O��l��V�hAω(�YR	~A��V��p�Xby�X���'8�/��T�~��my�T��_0�ߢ)Ga������6���=�?O�9x���
�b���;	��\�F9�Y��C^�7�P��\#�g*��y�[k��ﶾD����4������@���y��-T0�9�ؾE90{Jh��.*!��f� v&��,��+� �Q�]�q�[��1��N�'�CGr��`Hpu/�%� ���]�A��I��7�S58��s�/	C��83��O�P\?������ҴY����H�83hu���FJ���R���;΁�
����<�A�g�[T��}Ѵ��&(�CsơAX ��Z_@K	qz	��0ǁ	�j��d���� ��j�>�l!+M�5.`����e�Ћϱm���{)�G�G���Y��jI'��|����0)�I={��=(��7��G n3p��Y+.��V�%�����>䖕��O���A��׉��6�O���AT���Q�� ��w�D����
����,�Ɂ���C3ͪ�O�O4�4|��4��{��^��;��u�d�D�/�!Z�
��Q׀6��c]7�`�0���i6�Wi&[������ԫ��r3�<+�W+Jx��]�F���Gڹ���#)b�}azW�xV>[���MH�\���#�O�f��$#�8i�I���7�����j�F���Va��S�E����}az�vڼ�\�A��B\!�����ꂻ�w�U�D1��I�%� dm�{Wj"ճ�B�t��47�m�-R�J��4�7&:�s���%x�pRz��P�Lg�84��l��W������j2YD��l�kQWn��/��R�}��H��M$$\��2�n��J	�Z���E9ċ�f�\�%Y�$[o-7����O�Eu�a1�����0D�� ^�\h�L�na���?��{C3���
O=���8J�2��U���3��v#q��S�@��R�����M������4w��3�P�&2ݫ(;�?�vYB�`Ԍ�YUz�R�V7����d����ʬ��K���1��9�cTp?�uFGV��yE-E��S�<f4�%��jIq~���om�����I�=O¬�$�	��0a>��t�� u�:3f�hv�iGSA[�U.�/�$
��K��95�zz������<����d1P�Do*�p�.�WP#G���0������.�/B���%�_Ǵʒ��dZlbO����]O�N��%\�!�[���������U��N��Ɏ��(c�1'!6��=�6�"T��?R��&Yu6��J����������G�r��cs�h^�eIr������*�����!,Gz��>�o�<�� ��n��H��'���!o����䗻'fmw ��.�2�<풻{Ӯ�T;)k'��kI��E�(�Ɋ��=ju��������T��x����<�ͩw�@��c~��T������٬�J-Ɍ}�P�D��s�r9Y7��3A�k�i�Al����9x	|���?pcڒ�嫛h�V���&�7�^p����9P[��"̦��8]����y�K��w�.\E
7􁃼:�|a�^A����M������
���T\�}�v��b�_�{O��W?
r�}EI�$�Ψg���ˢ���{J� ��&۽]S�A��S�	�u�yJ�����,	����8"3����+���IFT���,�U�E�d�Wth!bZ	���e_O�M���5zf�V_��T�i�̶(��?�m��3��{�7��͇����a���!T3� 
Ո��N�g�N�s��~#ՈO���f퍨���mୱL���]5�d�%��+�j5�[�٩�#�{��G�=Ǎy_�\�r7_���s�b
{���G���Ke�;г�C}1���%��� ��eVv5{{eA���CP��
�r*t���ı ���`٩� ��u��G+|*�M�-��x���{�8fJm�jj�L/ą"L��L���9��H)ɥ�?�(�~�}=����vZ�>S��r�)�k<�oi4Auu���ͧ�����{E���f½�����c�S�?!����@���L ͖G�G~�V'��F�V��
�)����V��.ݠ�J�����ς�U5ȼ�؋�6wս3��̢U�z�tK"��
�<f0f���ˢ��d��)A��8������ݒDz�B���H���x_�V
5sZ @�+VD�@�|��u�#��䜲E?b~f���.$��v�$���������@Q�	6+RsrS��5b���"��n'U�lu�?�}�FĆS4c��H �����a��dqbs!�,�0��y������|a�Iъ�!ǭ}�<\��]���5�Lo���"?�>��9v;�=|=J�F�q���mE��,��0��vc����l�f_U	�kz�BH����|$$8/x��.�@�[k$��u��7�K��e������Yki��?*Fl�,Y�;e �����d�q��Vc��}��w��t�O���gN�ڽ�$�FьȂI
��/�'5�d:^Ts�<��Tڵ���A%�tR4=�$\b͘xb�\j��:�����6..#),�+We���5B��9��#JJ���]����R����NcFm̦�޲�jЎ�\R�v�<	ϱ����LoJg���|Q���N%�w�?���ʡ*�&I ��<{3nG��J���nx��~[�7Vh5<�J�,P�ѵ��ˍ��ܲt�y�
�I�暙�^K��ť(�k5�yMU+����{�	��	��)�$����O����$M�,���"c�a�|kq.B�v���"Ҳ���J���v[|:�uy�KIm>n9�LikE�`͠��Nҭ��5���2
w���(��mLvj��8����C��YN��2l�L1'�8�DF"`��S)��t2��ck�{�m�tey\+�O55�BqZs�����-��q/b$�G�ƞU~��2�������2�\*��9��/�T���o Fp�����?Ʊ�m��ĲZ���{�
C���?Z�(�����>�V���Õ��ؚMj*�SR���#Ï)�uC�l�6��s��˱�,��0>��d�h�sO��2�K[ncα{I�m{�g�d���-�lE�P���S;<�ު-�)��e�t�yMH]��	�)E�<�����q̂�|h;�����
jW5��٬,�������+h^��Iˤ4F8̐��/�m�?��8X�,��4@*H���W�A?B@L:jT/�Ea��f$hU�p]�ͩTW�8*bxf~/|0{���/�79���I�@�l�l3Ol׌�o(������G����OMC(���G< �vKG��ҵ�oK>9�������aлڟO�$���Aۤ�E�d�Y�G����t� ��Z�<ΖS�h��ْ�'�܉�ۘfEF�(�M�1z�X�Jɺ8������y������w�z����&�\gj�/K���]1�ЮqIP<�ǜZ�	o�²�_����c|�хQ,�c]��01WCf^%Ri�,�{=����878js�F�@ۣ�x-����ԔQj��y�-,�KM�+a�:�ͅ�W�q*8��N!&�H���x�f��@V���5dR���,s]��e���ft�]<�Dr�6��d�ǥ����+�gnw�孲y%AW�v�%�UR.7�{�3���^9 �?pT���c��/�m�\qrv�&��a�c�c�a��l��_�ԓѽ��\�����/h?��"E���u���õK[QwL;X:�؇���S�j�����>�e�e��n�|�.@�dS:7���µ�?��q\�dV���{nY���Tݝ��w�C�|������V�:�Y��YH���ٝ[A���)v!�2YB׉F�bH	F�?F:�Aθ*/���ϟ.B�m��;CiIG�L��?��b����U��0�S]v�<�f/�!z"���T�~�j;/'�����|�=� �;��߱*e]ɥ�a�D�Gw���2��ކ3�e�nEԬnI��ş������EAS`�g$���lȫ�$�@S�8�s�����F�دK�fn-RQ��ϧ�))Iҹ���)���fb]JX?�;���[��iX�<�@�q�}�x�OW,k��V�U��A6�"x��3F�����xk͵��\v
6��|Tl�;
���=q�6Ag������d�l��2@����K�q`�$�����J��;;�Nߤy2�,E=P���E.��z��0�	�J7�e�:������n������y�V��_�Y�y1Sd�Y|R9�R��e�һ���X7�ׅRtD�7z҂p�M�$�rD�[�P���|2���p�5�
������ՙ�R'������T��h RkP���R���w#���n'-�L ���cW<`�#�p�e �#+���w��fY����"��mB̶?��oGP�L�k�풿[�4;�x��Ap��в��!�'ϧ%E���kD�U;��r�2��Ѐ+���O�a���m,�m��5/�EgKϘ ��J� ���'� 4@�Q�@��,����Ⱥ�/{@�mY�=:|Y��u�����FݒS���70���ep�f"D�f��S�p�$&�U|�a�G���a�r2G�?���=*[4�U�p<H�RPp��t��&g��q��oB�����i˻�9�(>�\��o��	����T3���@%]o�Ac�%���ɏF��� �2��*�6��X�Ci��`Ŀc�(��P!Ѿ�L�?(f���2ax�ܰ~M�(�Ψ ������ ?��/�C�бv��[�� y䣩����{���@���Pt�XX���:�(��m���Y�̭|$��zHh9�M`u;.x�(���X�y����(,e1{u"|��#<����5V�?z��@��b�[�E�K��!�1�US��E�#�r����9�߂b�9$Gq�1Sa�N��O)�pgw��#Y6�C�JNLɼ!5݄m�<��Ī���*�񉳧��"��4:�i� �0�i�i%&����^��$�)Wu�S��;>�'��J�M�U��4ji�(5N�O�$��q"/���34O�E���㴇����jto+�6�+�,ŧCoC�N�LV�<�w�a�@֍��!�ݳg4��l�:1N+��ڟ�i�v��;SZBJ	�W�Gx��	��*��Riq�UںyT{<_r/�Uz�N� C�|I`Q���o�D���]D1X�~N{�T-[����Z�ü�\�ԩ������\W��Tf	If�#ӕOT�I�n����M�W�1u3h�P���]32�׽��H���J��驴�>����.��i��c�zk0��=����/ˮY�]��pX0�i�j�n���h�H:�nFF��'����ZV�ī�����b���tP���,�'�ƈ%4w���E!�M	XQh��0��C�)�9$��D�o[�N��Zt�h�3Xp��]�O�(��N��)\����h;H|�xcG��jΝ�X��BP��s�qP�[����xƪ��7�!��Qc��v��E�ď�j��y3Β����ZD3k7k���:�i;r\����7�RW��a��)�~���*b����
�Q!����Ճm}���癌Dt�ݢi=��*����zP�V���8����2O�-�����"Kr����Nk�p�4���n��l�(i�*�ڤ�Ek��_�
H�s�S�R�)%��g�v��UBRY�w%Q�w�����ǎ@�{oqr3�q�����J�����(��_��o�k�Zd����� ��5S@����M�%��V⚪��0��ey�i�*��ܦpj��<��a�`��|`PB�}�5�|��J���i¨(%(����Oi����=SʰN�T������������������ԟu� �WYm��PVĿ�)������w|��ҋ��DAw�Fo����9�n�iG��˼2 B�QP�i�~�0��� �xL�,Tpgm���T3��"ӡ�M��C4�h��ܳO�O �^�$����ȑAc����n�!g�Ĭ�k���g����a��Sק 9�*��i�a�g`����j�)�Ee����@x�m*���lB~� �@�Sh!���#1�eׅ-�m�(ޏ����[�˕��IF�����ҫ 8���f7��`M#�>1�t�P��Sf��1���nY�\8�N����V�鳩��;X�?s]샢�s�1sapbь.�n��M�i��m@�����p�en[����s��|Mw�C[8�T���ZwxE|SLΨ�'k�׵tQ�u����Lu6�x�fY&���^���җt�	\A��g?8a�R�Pe����P2D�s���:��iM�7��<���2���"I��y?pUХ�g��j��m��J�}�:[�)2�&��[ė�!�a�XT\+%��<}�Z}R%�"�5���[��a葦�S�u�ai#`\J�����A1�+�#\v���Bl����y�Mvs;��ie���� ��|�W/�7r�8Ũ��Q��0i\�m�����O)ٟ����Պ(��g�&vy��z��N�=�?&`��@l�qs��	���O�=l"�t�K"���Hv���iKU1�8�ץD^H�����Y�f�ZÍ2%|�o�k,(A���R�wFȰj��iGe��(�����Un��F�,�E�e�:x����d��Vx�
_4���!��4���h��6-�B'���]��N���D�1ͳ��t3G�5�E/ɿW��U`�0G�s!��E�H�R	���YvЃ�&.#��޾�u�;���"�ԧ��G���8r?ȸֱG�	��>A#l/�s0 �l��=��?Ӂd�Q..!21�@� ���\�N���!��iQ�)Z��K�*#p�}>09j<`J�������zp(�D�נ���mi/|#�C<'L	�[���n�� ��y�{h���\hNz9��X҃=+�_#L>{�6���l4��P)��z��l��Y��.�XR.��TNJeWQ.�����r��'f�@�Ë�t;��VZ��:'���-o)bl��"^�8 �;[Y78�0<�o�M�Yd䰤�	�J8�m�ҙ���c��+��	|�i�c~#�6o�i�-��}���_;k�9,�Nu��U�R?�j�%���a�)��<v|����{�$CO�3�Cn����,��������o��m3�i�v��z�O��f�@w������ی���:����0��=�.�o�}�rO-�R�F����e�L���8�H����AX��L�&��am����l�Fp�.�eXC�\ZR;%_~�5,}N����s�ݳɕu����X~��Ƒ$V@K뾼�8�'��q�l�%ۥ�I��U髬[��"jS���P��K6�D�C��w�0�YY���A's��M�/'�<�p<J�-�x�+V\l4ڊG���㦒ᵉ''��gp�1�JPN��
�5��~W[���}�,8{�q��o��8�}�IX��|O�WD��p�"�0��	������~PNMBWtM���9�Y��]�O���s�E���q���z#g��M �F>Ȁ-���>{.c;�$���a�}�xaU���������e��y����¬�~�����NS�kc���DI��#ߏj�s�-��ͦ�&ڷ7������=U��ǃf�f>����:�u�s�l�!P�u�#�6vf���0���/�Ii��D~���֌	��p`����B�����i� �-ˑB���>zK�w��{b��E���f���L77 v56ɋ�BH�X�c�DI�p�9A����e�g����a���cq.���P��MV����R�(y_#��^)�g�D"3���d���ډe�]�^S�c�*�������8�i���!�����]�8��o�H��8����s�<��jq`C���{�_�N�S�����a�ŗ��{}a.j6����
=L��w!����ݎ��gOu8v/��֏.��""K*����������wG�t��Vzs��ň���<�>S؇�Q4<�'`Cba6>^.g�X��4S�}�u�gBKb+���6��P:*f!3��W&q�I<��8�E�9A"���Kz���܀���&$sH��v��豣W� �� �5���u4RP��+�;s�	��xeD�Y���HQ��������v�w��.@��=_^ENO0xL����!8J��A$���ִ�%HT�^$������\=p'[1����K��=L,}^��y��A/ ���ĥ�B5��*9�c��F�-lO㴿��g�@mU��˵���	z@}}�hZO�w�~�xw�,��p]�;PN%WD`����������o�E��ݙ���0�?	W��=��o�x�V$�Dcތ� [peGa�/ +�E�]��w�88�},6� ���iq�<AL������\۫�g���v�m4�=�&|w��_AԷ�m�T�l������P�Nkʡ=�}Ǟy���Dn�et��^����o�U�B��bAy:"kT��F]���J_�i��M�It�t~K���}h���A��0}l�aEX� �	��.�
g�;�a�<�ژM�ݜ����TM���w<��$��	�6��y��T9u�	�C��x�W��w <!Z2ŕ���p�{�=é�C%w�p�!��Ǟq�R�������9z���`+1���#bT��
�3�d�2c�()ě��/�{����u����1s^/�;Z
�C���L�6��h�Dm�A�eɚ͕2sR^ iS�PՅϤ��jlFL;���LR����N��c��
͊��gPl���;�E#ͷ볏�f;����p��b�m<Bp?�Li~^=��:�9�)���9O��o��/�Ҝ
�D�*�Ѷ��J��P���5�z��,��~�܈��Ce�*w��L(e��XpU����;�)�kR1�&eq�+�~-�b���E�8�����cJ�ݼ��q4�u��/P�)CH��Jo/4��Ð�\˃y�6���OE�"A�<�ӥ�����D��}͝<�����	�P��~b���W0�Pv�"��q��M{��Ǳ��)rf���MH���ɀ�1��ZN���j�<�{ol&f<IE �5oP�:[n�~�~Q���J��u�լb(���ۊHaN����{KB�(��8�A�e��+�b�ǏŊ�O���?X����е�ח��4I�[�0Z����gpb�+a�7Q,��Е�.8�~If�,C��{0-��# ��j8�K>�Ҫ��?�snA�_�;�y_����&�M��������b���9���#�9 ����%yC�I����ܣ�����>��������T=�{���h*�x�@�H�s���$��V�@���-YҨVz��rV�I,���_�p��1�D�y���"�cχ���l��>�s<ԗ9�X[��&�x����G�
�=��-��)<��eN��BX+O��:�|R}���Gg����Z��ku5~���2`b���Z��A��0��y.��X�d˟��G�ZW��>D�q�x�����	��Dp��������z�`��+6(����]�a_���
{��$=���E�t��BƩ�a}��2�!���9-�xP)	�e�QuH?���G#�	����:۠14$09���Q.,BG��ģ+ғ���2?5ф}��Y�K�j �yq���P��%U;1���B���>J�ǚ����c4�ߘ3r%̑@�S�0�L�%�0�x7��Egl�e_���8���y;��.�:Z1�{�"��)"W����0{�h�����~N���*�MI"4e�:�꠸����s-9�F���p[]�}(���Y�%��>��z$�QV�@MƷV0O6v���Pm �+C��l	�媲ySr�Ҁ�zE51�Б�<υ3�bP/���Sx���(�c3�����3���%�Nu��]a�<j��{]�~�	��e���º?�QcQzx}�R��P0*�P`]P�*)��Y��r��� t׭�`@(�q�֟�u]���ޘ��Sd�s�b���_��9ֽn��K�|�㨯9�ևa�ĥ�O$��$�����F�d����d�<�3v_*Y;�HjL�p��H����Y�`�j4st��W6!��\2��{�D�=�Q�Y �D6��!���<�?��5<�*��\	�>Ĉ=4���|�Ә���%s�]a��N�;F�Hm��q+���$����@"��|l�j!�23�̻���^\��_����CՉ�d��	���O���$?.���3��׻Cڍ^�Ӫ�oN����pCQU��##u��܅��.[�1��1y�.y�AHN��9�z��4^�D�zX�EX���m���T�6)ūqy5����8\/�=k5-��´r���'��+7����.~
�q]y��{�V��31���D���~���|���i��wT7��'�0	#�z�`�:@ȀB�oXN��=���-�2j��`1�`bR�ր���u�k���.�/���Vu���'���s���g�3?ƭ�'��J��&X�X��lS��%�ZPO��ZﰁX��4��̜�����6 �l�z8wI�=�3�N�2��1'�y�l�'z�at�ϳ6����n,[CM~ղ�Z�k�7�w��#l	�ќ���4��1E����e�1mW�G5�Kn͍>T򳯍z	Ik���~o�0_�q�!yAM,�y�]�>b 7���/��;	!y�A�3��Mp;�'5D<,�D*�~dz��~�PS�|?n���m}b�u;��j�N��(�eX���a��^���v�/v�e%x;%���v��~��T�k.'�����++��4�"律gX�I���M곃���Z��5�L�A���K�~�:��#��-~J+��Cʭb��P]�- ��\)ᡢ����/�+vղT쇞]>D�?�P��"��d��̮	(rҦ�A�T>`=����2YS�^A��\5�,2D&�9���\jM+��,LM�(M��j���%�P�h���,}�a<j��m�|�b��7�9QG���	!�wt����X��)��E�O�w�`���S(ǡ�hz
�)ܳ��6���s''MV{�/�~�ʹ!Ç4��O�Y������+�A.�㰐$k���f�L�}i���K�<$��\�L˓��1���i�oju#�$��SN�ƌ�2g���Ɣ4���c��3�ܑ��4�ѝ��C3,���6M�"y��{�"�
��)� �]/j��1cH$5 �1�\R�δ~�>���'nQĜJ�$�f���^|���۝��چĂŉ��s݌�%g��t>@�Y�.��(y��;T�E�V�Ƞ���Ve����*�#+�~�����E(8��G��<�s�{�G^8<Yc��M�GQ�g)�)b���P
��H �C�+̊��Y�#Ov<B(9Se;�[�,����6��j���_��|���5y��UQ����F��{�~�s��>r��2\��RJ��@Ms���bK?:��$�-b�o�ս����JqI���'�J&ђ�MN��#W�-w<�3�h�^5{ ���l�X��UX��Y!����uaW����pXd#���v�3�SѲ���µ�3�U�`}�/惆#��R�Ѷ��%�Ա<1V豈'��d<�<' 8�`Jo0��t	�9�Z�Yj��eà T��9R�a����xÄW�E��K���fxGޱ��{l�b��Y�'����,Ҽ=$����q�����j��̼q�jnJ�|�ˎ	5�
����R����P��?i]/�p����W�W����H�7��qk�H�b�ug������gw�j4���<�p��6�M��g9I<M��Q�w��
�1Ǧͭ�Q�8�^��c�?vC��.�� �+���W4ߍ�x�p-n���K`�����'o�j$_+�C��z ��Ee�ѺJa���S8��׈�HPb�-B�G�O�Jz!P����s��ɻ@��n�M�E���\�)_�T>��ʅu���G�!�{;�.&��d�����'r��+�<����8�G�Ac�t�Ý�*�qqw�挥��T�%�n�� �#�s��: q9��~�r��7|~���H�뉋��`�����zrG�-B㥟c& ��x`�1ݢ� �ߖ���\������	K���.�ڌ�2��F�7�^�֓����|������Z/�G �b�h���5Շ@ [)�g����q�</x:޷Φ�%�a�-�t�H����~���~�h�N	7;І+Gj	Y�N���+���$��;�6�;w�Ug�b6%} �c�B#ǒ˷4��ۓ;�q����FEZ�t�䃔����N�S��_$��������x�n�f>e%�(�m����eF.���7�}J����\�mAZ�:�.b���;���s����
��@!q��@4��B�Ȁ�S�ٯ�k<|3ӉD� 	O����q��������@� �8h�dR<�dף�.�a-��x_fK,Mx1�gL1���YE���qθw��)^�-3'��ÄJsX���U<w�Lf\�~��;N��ɓ7e_�'�����,=�Y7�=`���}��ҙ�J�w:��C�FP��m賯A�g����D�H�D���H7�^=e���uY��Ɲ0�Y��z�7i�J 5��SЙ6��P�����H�G�=8Z�E��x�0����
f�R�?2#���z�+�V_���f�±���#=0eZA��m�\�t��e+S���I@Ԑ4���R�ъ��=s�-P�)W�-�X�KS�D����_z�Ξ���7�t�j�����Υ�gB�c���b )�\ʰZ�Þ��2�ر��ӈ 0��ў�1��ژ0?B���,7������4r$��^�8e<�`k
�\�S�Sk�4�E�b::6p�����)���~�I���񕕋dB���.J�櫃���k���/]��2C�nCE�XN���_Q�4���nlDu@�JX���~��''1�x`��*{�PyGu�v1	����6���Q�5*�9�~�H�S��Ǳ�;s�5~��"��ԭ�^6��i�c��`?g�Iܦ�b۬����$� ��s�i�
�ܻJʑ��5XDg��		��Ճ�2�>���:11��P�)A4�(�.�\z��7����_��<�R�XK��Rb��qRe�Z��N�`鯄 ��|���նibh��4���az�_�O�hQx�s$�	���[T�!�[�\\��D��G�3\�x7��~�lfv����Ԯ�#���x��ɝ���mb�@y~:��e�Ёb��0��P�ȦZh��Nv���<u��E�A�{���n�f�;]0��Y��L�MP�4����8��ڀ�
۩:�����L*"YW��*�?�]��x�a��ү�l�"qM<G[�֏:u�W�a��Q���A�aIZ��/(��;��4� ]�i�d��!��,�mvf 9���N�!�2j�+��e��!���C.����Z饬[�J�w��KN$M�
M�́��1�#�*�L��J���Kp�rd\��h�5�D��\�o�@��H�T5O}���0�9��V>EԲ�Y	���pCt��P3�L�l��W�x<���=�����*3�yz��==���&#�2�w��n�X�b���"龽��,
�4ĕ�~h�!���%b��RC��<3U�>�\�S�i�lA���l�C�6���/*�]�G��I&�<���7�םD��l%��u=c���e�%�%�(�	���$!x� B����s��h_c���d1������|��# Ӡ�	~�\���,�H�ň$���W�H_|m�������j�:Hl�c��z���߾_�o�Ϡ˵բ[S-��0b��?w����ޜ�`'D�a��}y�%Է5��J�?:A��ZzB��4f�!N���)���Q����ns�.0?H�n*�i~�錫�G�TN�<L�D�^��LxS,�Tʣ�u��2,�: ���pħڴ�YEc)<�קp���[��^51.�x��9���UU��`��e1f����׀�rAb�[m�_߄�@Nq$�UxA��LȲ�:�"4D/w��6-�X�SDV�� ���%F�E!�Kw��1��$%��ܹ).�uN�Ac��5�&��S��0(aj=���A��]��Hg�������������x�MJ�������rgOM��=��������y��4@�Qd"K3;�0�%ә�,/�o'{�S�@u��� ' �Nq�"{8kX����S��] �}0�?�Y}���3K�@fϣ;Hz��]�js�kIO4FG� +OD2.��'g�?$諄(I^�l�+r+ʏj�:Ye�KRᮢ/�?Zc_~�`�u�8K6Ӊ�d����D�0��:*�^���w�q�(͘�̟�D*
7�o$�ߐ�~���_�T���*Z�Y�<��W7���*�,�l�&l(����=HP4��#s،�©J��Vi��k7�3��h��3�М<��V[t�� �#�H�GH���5q�L��XUA1��jӺp�/��z`��u�o	���>Y";�ls�h��������ßU�$��>�Vx�T���IY~�L㮈�k����n����jX�1ǡE�&��rދ���^������-)�d_x���3PC���W��u}Z��o[�+v�p?�ϐ14�b���%A�Y<��*B6~Ο`�B:30���ԫ�%����ي�.+>�	�����j��@-ֲ�W+7��W�� Gb�V��/��(���Ͼ'���#�в��w���j���N���	�q���y�U7-x���~�rs��!��WY�5W�f\#��0��ޢ�X���*E��S[\e�y������&t6;ċu���W�P��@mS{�j���24O ��	��hE���D	-Ȓ��zF�
R=YxFJ�=�gܦb#��B�߬{|�+鈆�١���:(�x�Y`�=��a#�d.��i���]�F��GB�0���D�ae*O�)_JF�b�W�����<�'�H�k��r�9L��~�l�[܊H�n�^�v+�h�_�����z����gf��z] �7�5�M��Ԁ��W$MK����S��lzb%��m�s�S�I�rx��zcep�k	��Y�i�<�|A0��r�G��ɬ�~*��/AD�F�����f��ǲqi]/�*-Py���t�f��ܫ��V���(��f���q�
��V_$\�[�=�D_����R|���	)�ZW��t�E E�9�^��(	4G?O5d�	���n�,j�Sm&�k�,7�Hɋo��w��@����=0�M�fF%��5��u��;+&��������iؿ���w���Y?�-�����*YoRg0�C��d���O��XGa+D�帞�ڀ�f����-@7l��kK�gR��Sw`����cV�P
-���1��$�Ƕf��d�Բ���'����v��������a��p���X��rp�9{+S#�v��5{aBi]�]ZB�w2h�0;Q[~�2����M}А�~�i�й��h���%���
�w��Ĺ}��H^3a�yU��������4��Vf��!�@����HFi>�a�Bm2n�B�Nϋ��E<�H�=�����B�4Xā��h�Y}�D�t+Z��@�(��w�^w����Bơ#\���GM� ���m��s����Fr�C�@�^��P��l$7�������ȩ�Y�0�b��ν�xJ��NÐ8��և�m�X��R~�`I�B�7)LA%�x��@}5tUb���j�̽������������)�D����B��Kh��z��֊1'�6�V�Y012�XK&j���`L�n,ʵË[adt�m�LYBZw��ڗn�&h���㇆�zE^�r�l}�"ؤ�������b�08��P�H6�e��8S������~Rv#�@�B�Qk�mb.��܁wB{��x�K|��냵-�K-.���YEP(�o���s���w�Ǌ��l����E�D{.�Pn"���,X��T̒����mb����l�����;~�s� ^j:�G1)'x3�}��x.0� 5��:`���H�C�0ڟ5����?������L�耤�i�6��	��(a~�舩Ҍl�YL-1�B���3�<v�Z�����e"�?+NI�ۺ�S��i\��U!�2�~�i�w����/-Ĝ)I���GsK��1�b�� V�m������W�J �	��\�z�~�Ta
�66J�CO���9�މ"�e�����mb0[�\7Ȗ?��������ߔ-u�ڇ��A�����A��J��b��7*{1&*O�m׏���m�4����"�?��4F\ޚk�:n�����kO:�w9�Uᓽʰ��*�3%XzNӡ?�e�NK�!���r*��#�.���h��A�FH�+6(7S�@ٰئK�d�3K�8a��Y<?����5�&���٬yHq /a�3F�7���ڕ}7o��tO��H�SGW�E}��*�l�h۬e��7O�C�g�XA�o�!^.�p��j��]�B�̪D�[�.E���8] ���pn8�-�0!+��Ö���<�(�H��UC3
[
ǌ;�K(��VS�LD�JD�rX_�l;߃��v�hdӰ�p��.ٙ����t!�Pf��d���q���r�˯���Mp�<����܍�~q>r�c "�j]K �
��-אv��[���#. ���P�k�Zު8�i}�!N(�����7|�݈&�J�� ��Mӛ���QJK��)O��@?ᣄ7�I�:0N�G���u,҉y�}�D�F��`���@�Q���E1�� ���1h�O��*�A�%�����k�M�er��E��:&�I����=x�g`�w���d���˶�at����n��Z=����������ͱ���D�D�������z[��*t_�jdƻ���Z1��{ ?@21b��T0}�,�C�XK��Lc���}=�޽JB��jr�d2�¾��<�g�1�<l��n����✕�Z�z�ɪۢ������b7��Vw��䍧.0l���k�L�H��zSC_%�1�9�%Q���[�OaDV�D�ⴖ0ke�� ���a/��4ڛ��5���nU���r��)�d��(`�V h�U��uS�)D��qU���'�bY_r� �y9�$oڪ�ht�ܹY�q�U���r�'�z}E͏勌���zG��e��Ȱ<����0�3�EֶEپ� йp��̴��c��Z��R)�Mh☝W\^�o#�uBPK��((�)�ct@�qwY�����j���^!n�W"��c��kS!��8���س�� %

��02J.�����$AZD;:�sp�A�ʿ�p��e�E9}i͹FvHm�$�;���q�m��������eT}�^jJ��A���	y�7^�W���H���n�+�#�V	��bE�'g���wG���U���l»L�6V7�,
S]����^v��R�J�>C);D�dp�0�J΄�vJQ����I���_��"�W��N7�'���� �{�7ra���+��Ѓ�8�?� ��;�c�H�~v�V'�I��S�gwi��!O�28���#�Q���@+.g�7z��2Z�������kg^�ݣ�6*Wn29����"RBH O|��X��a̹JsD~Z�}I�$@�+w���wG�����\ۋd)cG�ϋ�P�����ʫ��;��0�w=@�5��������{�%���FF��ǉ�~�χ�����~�rw�)�-�zuAi�c��E�c��ԣ�x{r�	��M�%�q��_l�|U��!l�t��^��@*�`���1���j߻�5D���[q���ui�����T���5�n��܀�ő��f#�R/ ^�c�(���%E-���p녳�ɨ�5��]!1��tt�cCI�"i;a�
�*��	�����<��h}�uj���>WVm�B�G�ҏ��'�E=�z��+�*�F{rS�wl��x�X���f���i�V�����bY|ĝ뉂�ɂ�3M
���Py.��V<(}��Z�E#>!�s�M�O�P�A������kxK�����Z����w��\����Ԑ�	V�A4.J���5o ��Y6���u��꘠x&��/�V@
�-.2�i�rC�n�ٙ�L�!��)P܅��k�Ksf�$mZö�eM �K!:��qgQQ<�}��a�P $��� |�v��G5R���/��jO�򏓨E+��7^x�@t�l�F�E�!}CF�(s��싉�~�^~�t��Ҳ�ymg�3��.�N���¼-b?A��r?4H�z�)�l|e�H��e�٘9���`�{�C�M�4f��zs^������^���
t��y�{
�}Ry��1w�گ�V��	�i6? 亙)+�KąB�SB!�[~I���dR�n�}�Sf�P�
:���Ρˠ8�a��2sJNm�8,(5����_�����%.i�y����ax7Z���l�G��Dz �:̬���y��h��@�q+���l`�����x����+d\��K��	W�z�N����&�o;��_�G�T���b�A���މD�n�h���;9l�KL��6�[��)*���zB�N3@m�R��%��#��\>J`kq�F�u�Z���نŰv$x_<"1�ݝ��D���×P:�2�!����P7�c���Ҭ�����������O�Ecx�Lx�����8�Ч	P�TN�T�������T*8X5��P����'��Dt,�A��sr������TN����F�,�F�=�
q𴙍I�=UH��Qc��(l�E�@��5$^i��LrX���s:5k� A��ԙf�&���kHj��.��'�@1l��}>��+P
��=�@��Z��1K��n9_Y"�*��D=}{Gxڎ��Y|\��[&`m��1�v�ǎ�C	���M�Z�W��ȍ�z�\����� άI�-�5�T�( U'��͈Ap'�Vs���0���Գ�˘V3����	�0�����ѷ��3\`ۍ��ߠ`�-��8�RmF2��:�Od�H��*�u�x��d��̻B���mm�@�D6��G	e	~fDuQv����g�5ǟj�H�2�D�"!�߾�Y��K2���f0���V�]�*�ǵ�)nF�]�
}���t�d��-��;{Dz"����J{����=�0S����FUsw�)�Dt��Y�Z�/�cp��9� �t�I� C�Hy�7Tp'��6��>�1PRK� (��P1����>_���Rg���^k���(��:�3N�Bo'']��V��}�G�l�jK�2�Ͻ�I�)Wyvz�C<<��kp8f
�����Y9{�a������W��" E�~�<z���UCY@��ҳct}K�gӛ,74m?f�.@|#�ܘ�.�W˵37�0��Hb��)Tv/��ǔ��ƝG�>W�K2��h��µF�~A^j���f�1+�ث�fcb��u�L��?�o�_�ITl�v���֮ȀF ���������	P$�Q��^i�]����}���]F����7/cn�J�ws	���4����m2͢�_��f�?�c'u��,I����;f�p4��_$N(��hNd�K�CXi-SOr��Q�t��A�A��=og��bbZ��S�ٌ����k�+t�����a�nN��h�}~$�o;=9�-Gl^�:	o�#5Ѡ��9�	Bs��vƜQ^���KJ}�J��k���M�� �]��8�쵦�+\ِ��Û�$�[���b�'0+�J	�GF8س�k�ͳ��P���&<�� XЍMa<W*��\�x�[j�������֍���T�s�^D��]Bvf�(�`q�J��f���V�������Վu����zB�sa]��n_��,Ɇ�u��5�9:��HK�Y�s�wF�߮��e��aj�^��|R�"�y�KB�A�Dd�ny�;q�F��X���)j��i�ޫ^�M
�t�4�7F<�d� T� �
Mw܍ь�ғ�i�_j�Zc���V�4jD��4�ֶ)���o��X�vC=H��@�M�Oq��$.�Qh��q������⼥Y��A��[�b�?Uv��Ij\�-O�o��6Y}��[+1��R�t�m�?,���tyg�Ifļ+%��{��0��bG��0\�u�CE��(�M��u�����Mݑ�p�-�F�]��I�n|	�.��Ҟl�M��ȍ����!�H$�9�p��)�k�����<e�ś�F����f�&���ڨ�!s��Y?������co��%a]DMef>�?�XQ�z��&�p������P�V$��G�g��8@C�T������A��]sֱ|�˳C���!-شH6�OO�l�&j���(hkx��~o#�=	�v"�Fshu� H1��jΕ�{4�4*�|����ܽN����a��<P�p6��cN�_i	y�!?����v�����}�T�b����B�yZ4���L|6���������O��4J�nG�ֱ�:�;�=�h GQ����j9u$��V QN��N�|B�q��ҚJ�%Q�J�b����gS��Ҩ1��5XDW���Y	���X�*+w�+��(E\�C���RU8H�g W8��՗|��](�Tps�鼲�myފo����SM�4 lh�۟S�9P+�i���:���oD}$z=/��E��#�䫂���v9OHy�V�� P��HFF9�Ӥ�� ���Q���2z6�Q�uh��R��Γ3r�����d����v,OSR	�u��z�RR��e��g�c�c	x�m�7�I=��L��D�*^����$Б[����{�+8����~��@�	9.�����VJ�?��i���)��f��ba"ք��1�SFg��Ii�N)m·�8�b��_�Z^kWJ���i�̟��Uh3EhQ�֘<��"��Y��3�cu�r���R�&!9�h�jⅺ������ڼ�ݶ��q�� }��ځ�d)��V̏��{��l��\�.�K�RO⼧�#�m�0�,��˝�� ;	��{��v����J����q��{��ͫM�	 �0"I���H�D~�m��CD�)�Ƶ���}}I<�g��J�C�.;.͙���t�,�p�c��L�:rj���3S��gb�z�iN��{�o��%���Ev���,�u��-�b�[[�5�!Ԃ3a�����^�b��>�e��V���h�	��λD�?̈O�6�ܙ#�H�d�=�1L���Ū(O��	�_�F��ܼ�,�ڊ!	��<��x��� Z����y�Ƹ�# w#�	�B7@��bҤT��EW�;��%���k(oJێ�e��e�z)� K[�S'Ʒ� ��|'D�x�)<A��OBp���X������I����_����p֯�=y�"�x�2<��,[:4��&b\v$�qG�6Gl`�O�`i��gzy�(t65����]L��ą���v+�c	���FŐ����j�ٟ�>`b��:�=�Mgs?�|����}ÆJv_�T�F;�+��激B�fVxU����L �2+W��2���h�b�2�
�@��ojS����!��A?A��V\�5�5qpn���)_���izG+Z���*ٿ�����p��P/<��}���3v �g�\L%�Z8�A9HaD�bG��"�ڊ!B�����w�DN}j�m���u��P5���$H��'ͧ~�Y�U�G����
$i��p����2'�_�7��)������,��U�8e�)�~U�Ӣ�����?�z����!H�����>���lMW����P�!�<�$6���7�)P� �*'H$?+�nt�5�_=F�b�ӫ�(�"�>sS}��x���^�
��(N�+b\I����"�,~*��6�E�=��^1�Q����$����]ʹ�FA5��mI�H aA^O�x���2�/�Q<��-:�+܉\Y�%��v>̌VQm���c�k�K�h ��#H=vt~��?�w���As�qz�5�%����뗝���?����QϏGJ;}qDܺ7f�Yq�5�'ֶC��=�&E�݋$� <��2�
P��8j���⠿����Ӣ�c��с���vY�l�5HivrGNm�k1F�G�c��g��ZϮԺ��o�P�jS�0wh��,���M���������=~������.�;b���\�^���w���y�O;������P<��/@��Q���"	��\j�`�][�M���f��R��j^Š�{��dP/��2�Z͘<+���4_��, Bq$�w��$V��D�z޷�;r��Y�� 3����Lv!���r�B�1���պ0�c�� �63"�Ac�ш�WZms;�GH:II�]I�yrLe�i��a���̏>|�M$e�DW��E%6�f	: �t����-�'l��E�d4:�f��hb�cH8��系�~^�3�����0� I���5�5~iI� *�L��j��g��8��Nɕٳ��Qn��~2���w�0n���vb�aigxe��	3��T����䅯'�/:���7��4$n���h�)N�f�/���|XE;G�-}�BC��x��d�4����	փ��'CO�>9&���"��糝�C3I��8��\�1bA�J��xp\���%�L,�~NG�Ho 	�e��kP�N���ؽq��8�6s���"���1�[Xښ������>Sv��F���=�00_t�U	��EP&�6�~t	������*�T����ʊ.��%��A��
��-�=�Ǒw��Po�g�NƦ0����ߑ�W�'ix�Y��$�\4����2�^?0�D�
�zY�����͞�ֈ��K|��8��(���w����EPJ���:���)(Ǖp��"�/w�~6c�1����J�>8�qk��f_7��[����#�����	�����mSk"&K$��N�b���Z)�e�e�Sg��Cd }q�ώP
+�G{Ҕ���CW� �S���PQ{�H��e���-�Ed��������f���(����;/�-Wf+�t!ǀ�[�lGb�|.'��IL�[��:Pt&B�~�4xż	T� cU��h"j����.�5���.l3@���P�
+u�bEO���v+��蔤���U<cBp��fD _�or��(���(�3aRI�t�p�_kgAR�>�?�ӈU�ep�ndY\����~��((qX���~���UI���|jkIr��"���
�P~���4�R��� ϩ��AӤ�H�K�����:��l�T��������t¸B(��s��-A��/=;`��>��J��< �^(p7&_f�	���{diU���k8DU��C���`v���* (���i��֜m��`�Ik���ӈC�j��4����5.��ĆǾ��* D,�2�^�F�|��r�t���b@���:̏�r�̞e��B���8X�� �#u����lA��^,��
$�z��aP��0uBy�/����Q��gxs%Tq{S�VuB��4Ni���HˀiN&�9Ͻ!�^'���`�u��ڻ7S��*���C��9qW%��;�؎��yD���B#�8I��yFRB�k��(�ĥJ�����ѕ;��o�s�34:�H�������*�a����Nb"��� �e��§�+��}�W<�
:O�j|�>�o�%���A�S��Mw�(x���sl 	]�M)"T��2�<�y��<6m��8WRG�������(bkJ9� ��jN���n�}iI���}\ࡏ�N�P��,{�� `��@"���y�8��.>'>>'��=`�;����������ZV	X�~�Ո"�_
��ǻL��_b~�[��D�H�c� [�X�I�b�e?{۾�ZY�̴��}��f�\��2����	�̹�=?C/�Q#����1ܛdA� ��s��v5�坷'h+f�dD��e�����J��r�NԸ�l�����R�m���G��:.�Z�9[ 9}b�p���j�><�|{\b�:J� �b�s��`%��i˽���F^Z$�rs�P�V��&ʵ�T�rm
��_.1��O
��-�������Ou�t 8|m${x��pX{�8Sg��+��6@�Px�s���qlS�0�KaNbx��r��,��F�$��j�sx���t�@�C*t�`ho3�|��l8[��*�f�5ټ��t'Q�pY\����M��X Z9�eEEFpᾃ\(ɴ��;�mY��^�A�E�c�*�R��A��?��l���$/�5@h�:^��:c�[1�&�ȧ0��?%;�2��Ū�re�[^�n=.�>$�F� ����������N�cCJ�a��@��O�y3���V�w���ּ]ޜo�������c��cj�o�֥`B���s�*�@k�F�A9�U#�P�mΛΆ�C���}pۀu6�U�r.�@��r(�䷹�25CN�0��&���21��Rq?�8>�	�S/��v~����T-��a�pxy�_S�H�/,�l� dS�PsΨ����C]�/��ay^f3T��՟�0l���|n�c�"�,� �Ȑ~����$��%���1Ȕc;��UcϦ6��/�H�c�R�=[�1��xZ�ʡ��JP���4%���$�E9�ç��3�S��u����QIw�t���*�lUn�;ŵ%�ۤ���	>M`=�|w|��I0�m���l��M	�o0���������*V�,�-bE��l���l�w��
%@��
AO��m���.΁�L�uP�J�v�|N1-"P��跞���]ie�f���q�<�.�RN=��IGD�f��Z��Ɔk̓g�r����:݅3���bq��������&#վ���D��߁�RC�X/MKn0-�
���Y�48�ϙ4�Չx�;�t�yCnٟ@b���x@�]�;�⁘�s��2=ꚓmʚ��n�bJ�Rr쓧ʍ5|��C=��X�T�CV{Iw{���`E�"�꽞E*�<�>��S��.b��_����@��1�H�\)"�R����5����(V%ҟz�	��J��}=4�dA��ڃ�]\��S�	j���q$d� �����>� ����^|	�Ѝ�>�i�S���G횐�����r��̳+(,]��O(%��Ptv(C#�a����W$�ؔ�~}*���;msj\�NuFpٸI��5��gJx�o�  n��;�nw&:c�e:Վo^A�]����X�l�������~keZ���+���ꀶ�����*��>a�آ� ��4-�/�PYB#�#�O���-����҂��}��d��h��gx�S�E�$s�, �G��Hvt�,�	 ���8���[���N����)����=?oH�#&>O��/Ň��&�f5��k3��� p�U��㏕� ��.���Oo��b@i��R�ҍ����	�z�u+�n��ҵ�t*~CE���`V�tg4��`mR�WH����%����L/�xO�Rͤ=e��_�|٬�Q-ic��X�,։p6o���o���!~J��Ԩ�r�g]�����,�+  q9ܒ�]�0e��2J�wV�˲i��tnK�~�߁�,��I��|Y=J�հF�u,�7�Ҹ6%��[�!*.�N���₦΂Z�rk�Ǭ�`�ɧ�0� ��ㄱ�y*q���'�DՃ����j��'��(��|�⽘��2M���1s0܌�7jv�O�[N �R�4�Lo��� h�C�34��G@��dI�⌬ખh��յA��Txn�=L�7-�4�xڒ�h�(ATOJ�Q���P)����r�Qp���f�e��������~%R~�,o�<Q�Ҙ^������:_J䢁���r�����_���Y ��[�sJ����+e>��귦���,B�Ǜ�F'�������+�A�쏳�Nm������9Eyrv���_�52!Bi�}�{�&��B����9�i]i��|��dQ�
X[�/��P���F��u�(��?L�yE���w~<�X�=:��$�}�\'��g�o�oN�����Oܠ��>��P7�J�
�ze2Q��:��$�Tkm�.A��nww�}��T<�������<��Mw��6��!%L�>�GD��2QB}���$�J�f,�KD�d>V����_NV�|v���`NI���W<q���`$���-�IU��ș0/f4��,b~�"᧊����$3�c`el����m^�K<�$�w*�������i�<P��e���C�Z��EL�jF�'90�&���*f�x#��Me,�f��J���`���%.�
�k"�r���;-�i�/?����c�u���h^i%��08�t:�]�hq�2w�R�ˡ�̉gj�B�G�uFS�xh_lW��^��f�X}��|�E�ؒơm����[EH-Ģ����O.�L�xH�Eګ~Ӗ$��2?��䗌Ӄ��BP�bB\R��wy���e��7�l�2��u��VCˊ6mz����Ͼ|�83�)N�-�$��H�2�O���X��RA�[`�������������7`���AmA���T�(������B��K;dp�	D����c�S\����S�� ��׆"��C$���ɂ�y=����ˈ7Ј{0}��$`%<��z|
�$���X(,��O��#�a^��8<C
�M�T^s�����"M�M�?M ���]V��H#���͝���"e��|��|�u֟f4��� ����z��OH�@'�l��f�e��k"{t��$ �«���5_CAR��C8���W�9nW����`��E�H���h.�R�g⹵T�E����~$�a�*v-�=#/ꩠi����T��P\�#�I�sM���K4��"���,�"�1�4SSg�a�t#�s��u�]��]i�����]9SPֆ�XS��cO�
�,d���ږ��#��#��̵�����1$������%�d�o��]SE^)�u
�G��髝�Q��~���h����9.��?@�P�fJ0�2��m�[%��5L�U�è�*Wx�օ�xR�'x̉�A������1�RS�diK��b�6����^b@G�!F��p���n��e^+�]ӌ��*�E�1��\P�b�0�ۥӁ+��iy�P x�9�a�"U�g�-��K������`}y�r����=Z��@ɸA��ɵ��q+}�Y.;�*N��)�_���y,�Z4�� _p��<�vAaj����	7X"��
a�m���������<t�}H��7%!����_5t�h�⭓W��j��oR�n�҂��M��;~!��B�a3�J5��������ϑ4�=�5�᱉�=��s¬H���˳Xh-����oh� �Qo>X?��	<����Z ���E5U]�y�/���%���Z�8�@| �B,K��`�͌SFl�H9��Wĉ�E#*�Y~��f��F\g�s�}����fy&̠�����W�N\��=;۶.]���/9�|�������;%F�X2�:�)�4�&w^��?u>�Z�Ls�΃��c!���rDr���D�ANÝō�MP�QyӵQI�Aa��6��[�E��8T��V���������웏S�Y��_dl��/S𹽺6fЌF��{";ϼb/���Up��y�V�kU��h�yiP�qr1����� �X���ϪRky�ɳw��ODɺ�oXC������^4�<q(0^p����f�������F��F��7��A������XEˌ�����)��r��&Q��%Q��k��<�0c��h���Ʃ3-�8 4a�c6�Ł<R�K7Q0�Ӳ��z�'����)��4.��Dҹ~��5���X���b�'C��X`7�~?��/��j]�+�\ �Y��U���p�h�������+a���od�*4iEh�8I|� ��N�@�I���ܺ�a�|���u���`�UF	�Tc<J���u��`-|M"S�y��V���\T]�hhԴ��%��?��v�5��U(�*q�xw
|W���q*�Zj����s4}&A&@�5K5�Δ��RS�I���S1#����h�3q�]���
����6����8��j��ATɀx\�0�[c	���eV�a�D��=85�A�������?��;�I�CU�N�����`���
I~}Zb��9��6��"����ّܔ���5�/����p��0߽D{w��dH�������Ҫ��Ӂ���l֥���������&�:���;3�KB3uG��d_��]]f�@���~Q��yuK����*l>��Vm$
6mkj�kLItmº����fF���3������0���n,�l;�.a�DK��wd��(��%��S��AB�%��")��J�3��,�֟W`���jRF���*e�P�Æ���w|l��^�Jυ�]d�/Xt2��"�.*<������#�c�lڸ|G|�-*��u�bg����2P�y����:ɖ��|Ӣn��K�P���arc�c%X����8/	W�ߜ��	z�~9e�����tΙ����։?�_��t��Fgh�L�Խ�.���Sv��4*�J �x�o�?��wc����A'&x�lh����r��AgX��4�6N��<���ȸ�	E{��9F,��x��-�,&v]n��x�qz�P}_-��>����3@�'��PZ�J�_��0?s���B��̍_�(n�g�b1dJ,� rYs��<����n�Nf?�g�U{�L�얅ј��	��q��gK�|�������I�*���7�;(ر��މ�}�I���R��M�)�ֿ>B)���_u��P���h�;M����[���k_w�M!.��[Alm�70Z�ά�lc�KU>��Vy�1�
"��1��5�U>��a_�l��V�%j��]�O����!�x�`�ZJ&E��*e��)~c-?�7 L��4o��:�':�|U�l�(�
1�m���8W%i�v����`�^���߭XX	�5�D�㰧x'�K�d��++Ҵ��.%�z�3�"cu��P����ڡ�L�"(T��\����-����԰��%�����[�^�J�Z���=^��&9Ŋ��\�N�?H_��SZID�l��r���-��a�i�H��#�O�	�X꓆md6^Ƭ|���4	Գ�2�O�ſ-��ǡ[�c�x�H��շ3A�GU��>ř�)�Pwy��r�22*+;dF��*ɐ��?�}�G3�	pޱ-�>yN��D�I6�-T�2u�Sp}6|�+Ѐ�v/)]O��vJ��.�o�P��a���>��g���*Zƽ�V��w�U-�>�i��v�z{��-��T���H[�<�!��i��F�&��yZxJ���J�\*�����=i�Z�M݌��8?�.;p�PB��ó����D9B�O��<��F���0�Qv� �k���S���YU�0C.siW�S�2E�
���݉�^���C-�[�� ~�CF!��v���P߁����y�L��<V�de�'@ ��q�H�ro�~��Xm�����Cp���YH��o�3
x����ϫ��i�+�$3�	��Ҳ�=�q"��v��&fM�)f��s���J9V#g��מ�3_"���>Y�˸� X ]�	��,	�ѐ��A�����-;�flBs����Z(;b��m��m�EH"�ZՈ�pbEV����
��$7��T($�<S��R`%-yVk?X(��j<"�Z��;QM�hD�����,��gnKA���\L���S���o��|�#4�E�\�As�'�2��X�Ϙ��y��&�K-�!Z(<��T��x�j0���U}b?7���hwU�(C�.c[#�ƭ���m7E߷�f���5$����Fa�kq���{A�,z��y�6�W�@}�,s���3	h�s��"r�:/�6]F��D��E��Wt��xy2�0[D1ptAy��/N� Dm�,n9['��ml^>
��F�O��lO,h��������^��Aɡ��X�z����ǣ9�Q�,����9�Yc��B������U�뽦���/6cCv�mNL�@�/ߞ�=0�f2����T�O�Yy��OuԸ$�P3���Mk�Q 6�1�;�2��fl����Lq��Mi/�{w0(&&4c7����7�O�B��s�)aQ���B��^4�}E��P+j��k��ȹ9�?��3�5 F$����T|����&i0�A�v`!vI�9|u�I�6ee��N����ajeY���?�	�&s�v�r��e�u�ac�S�_|}���s:3�-4�&�|���s�hē���0�,1"j�!���ǚ��GOj�=��r�z ��%��6P����,�l�@:o���_��d@�ږJ�Z������8�ÅQY�[��#�]��y��������J��gjw`�jO���ځ��
Tn?�	�4(�����~�kLPm�g���p�i���ó���s�Mc�r/�y�xg-�Q�G8����d��0�w'5��Xb��$�K4Mjˣf�0�P��V�Ë8�>��	~ĝ��e��<�o�Ww�p]�-bɅQEY�Ҷ�!v,��Ef��
�RڛbN��o��F>�X-$��Or�qq�=�rp4{��|�M21�I�B ����t)�Ƣ�Fݡ<�{�w��=�L~�5336���S��aLF�J �}W�M�L�K����Ȯ�reU���+��g9�	���6�`�z"��tX�W0ǬA#+��t�$c /N�!K�iډ����/���/@a\Z%�'^dR<ҳ�@3b�BY*X]$ܯ�K���k	ჯ�qx.�b-1p\ʸ'�x�e]E��@_�I׷���y3�U�ѷ�^+� eBՖkz�eMz�#(�<vw���o����́�Ƣʵ-�pAX�X���3�		 �9����58�D�6O(Wwj&gqs��4(,�/J���#S�O�J�)^:en=!*E0�ժ·�N�8���Ʒ��&�:%�^�b �v-�t!D���^)�n�6]ep�6ڋ�ϥ���)�>�Q������T�JY��k�o�lQ�l@|
����.�CrK7�9lK��n��e�B:䲖�1�d�n������}���4I�v�̝�J��%���+�6(�k��ѿ���t:8��J.��C��V�~�Y��V�|�3]/��Sp���"L0B����&��C�÷��V��¶�=\���{���G�+�[+�j��	V0���?�<O��0%��e$���l�%��G��L���SXB6���XKm�!�=�o�Av�����-�=\�U$�NSk��K�*B�$�IV���(���Hb:�[d�b����/��u�C�ܪ��P?n*މ.zS�Ǆ�iH�N���9��E�Zǜ&��!i�H���I�����c����@
\`1�7�6+��q)��_K4ceAԛzܱ� :�4��ٖ_��%�,�zި�U�sP-x"�	�k�<=.��~�-]����/f__�[S�@�q����Oe����W9Ϥ!>�?���S�t�,�~��p�I��⟱��Ň��a�8�2������S��?�u��_�J]�n(�$X��َ�f��r(V"�F�C�c?^��w@��4�G����)*㫰#n�J� ��^{(���X�H���DX(��ӭ(�p������b�h;��r�;B5.����|a~'A��~����kj�5���Xr8��'Ca�W�� P��h�O��^� �a�\���U�/���ѿV��q�4��*��M�&�����C�v���|3zYP*44.������-�:��YF�3	>HA�4F
T�/�pT��r�R�g�ź�eΠ<�
Y�Ol�P��=U�E�}Q�F\o��Bk��3w����a�6?�{ՙ��7�����]�l*�	R�^4=��],�L�.j�XY���'[X��,�[9�V�"b��m�������6�l$�㛜��S�qw���|U��:DSCl��@��ũ����#-�}��5�=���G��q��o���`�8BN�)O5��c��p�f؃�b>��Y�����K�q1T���5�N�����KA�I��]�H�q��uQ_n ���s�{��cfXff�9sI_�#B�� ~1����W�1��v�FG0�/�}!�p�䃙O���A	�y]�s\���z,����8�llE+���7�Jnz�r."a�J����NA�k��i�b��Sס�Y�|�x+��U��'�B������1�U`�g�Gr0[��"ՒIF!��ϥ<�����y��k�O�?��6�F��i�5	겟oB·o�~m���s;�l�P�E�b$�:�������om�k	ͼ���vSz�E�$�v�AFg���&Ǧ\u��f�S�,�Udj�;����7�M�eM�C�^���#F� ��=��K���y���4��13�9���PAc6������D#ƍ�@�Yq�ZֶV3�Y|��&��1P�M��X>��w��w�L��� �eq�m���믶xx=��=����a�*���&��lsB�+D�Q1��V1֣��Ń��q.MZ���8*����Z��Җk��c�����ͽ�e��]ȭ]�:�ؙ^��'`�N��W(�Jd{��E��\r�[w����h��_�H�ȹ��!�;���~������'�=?���A�q�ՙQ����9`��jt�/Z41�F/��M�=�mݑsc����0L&S?�φH&�.G�������.��W'�t����]o��zƯ6)A{<�W�*���6W�Ɖ��7+�)�,U�!�7Û3.�������m���vY�� ����/Y��=�4wOF�Y�3��ʦ�w�a�T\!����m��	�P����W�D��h���B� ���b���2��^��=R1
��>xj��5�t�}�=��#"�X�%Gl0)��Z�1).(���7�8r�q�ZU�J�e����B��KT{��k'���ק�h��H�Pb��;2m���ϰB<}UFҳZ�!x�v\��w�l=Ш`2�}H�Ĩ�� v-�0;�&��E����a��/C�PUȃ�?��j�a����F�X�q����n0E�F��|��f5`Q!/���Y<��mp=x6T�`�B��{䔂D�M*&�)����!�洨�@�?���q.���X�[�L�򚎳)�C`�Zu1S�r��,��.�ޯ�c��/����U�'����|�k�����A��w��&c��o���j�|3|$�#��%a�}{8u��=Bt�Á{߯��en������YZ��n����4C�DR����46���&I�T"T�Gڙ�G�i�������bT�&��N�e���".��x	J�Mb���)'��^����}�vjȡ�w��A��/��׬��#�J�yZ_�q�7l���@'��֮Y���dk/W,ye��a��؂йn����7@_�_4�K ��ep��ӸIN�^;A8��W�/'�ޑE
���w�!��Br"��p��O�!5�g?ۓį��]�gd����������I����{3j���>�Y9�nJu��`a�(�F�T�*,d����
l�X��~_�o^�C"6"����:Q8T���2����S���ǔć���6�b茑���p³L��X�I����F�Ȗ9<�,��4)��T~9�`�����r�'!ȃƬ�_�s�N��%T�A�ך'RuYi�Y*f��9�q0A+��^�陋�$`�W[���L�W�p;D��{�@���t�N�Ӑbm�U�]e~K'�lw(+� Ғ:2,RJJ t>-��#@���9ЎK�� ���Ň�,�Ư�:�z��u�:ۮ�fDr��x!z`���^��L(�.�I�}q�X9�m�!Wb8F��:8WX���n�+�$+���eȱ�n��ݽ����.`�¼ء��%XQ��&%0Q�y4o��-l�`R[g�[Ӌ���̗�&�G�4�%�+N{��J`h7!A+R��=<G��m��ƍ�q�����0���L����U�d����^QV��"p�����2!]$�J���J��3oB�ް�,it��t���}����SMI���N�XZ|�|�C�[��x�&�O|c��I����y�+hZMUnrAsTHo��覯ˏ��C����ώ�ʻ�8���]��6������?�!�M�CƂ%Y��Co:�[�Q�k�L�9����B��&�b���`�iS����uU��#�RLkX+�-v�K^r^a�T�>+ր��G~���x�1�
w&�V@B5<�	�|RQg��?�;�-�φ�D��PH�.�Q���2���}Lx�Kx��A��9�W��NCW�2F���B��;~� |�нֿ�c?���͐�Y�;�����y�����Mt��o��Y������Rh*��LyJIx`X�&ζ��Nt�/{$�a�@��P.K[�.�f�j���$�����z�E�E� ,�z=7���H�)ڃ�uR��x�5Z�� |2Ґ$�/��{�[5	�+Yۯ\�d~�^8Ƀ�gO��������]�//=4�_��6-7�G0d�
�a��5�5�p��>.L��/��zs��*0Fr��2I$��tV�%X@.NV>rd���.ӫ�����!UPz?o�؁��[GmnK�����\S�/q����`�ײ�Q5怺�C�23��,H��+J�`�r�u���*ݰ�=�2CFl�#��8άډ��֎����p8l^XJ�H5�������~S�	�F�i���K�o��$�m�U��l��be�G�g<����I-=�o�o.t0��$�ؙ�F[�n��2�H`�n����<�u��y��q����]
�,:?��N�*o%g)��4�;�}��35Qzު)s\벤�ͨ��H(��J'o��]���'S?~��3
��1Jqz�g{�c�7�UbZvz<v�y+ �P��/��Y坼 ��2��*��c+]�a9H��}ƪ��J
��%�䋂��Cєjrt.1֦$6�r��ʊ�{F��3
�7���ֹ����[1HV�6�N�̀���w��oA�y��%��3��������o����c?�7��	VX�UԱzBN}y��QZ�hϐW5[�ς	逽t��{b�AF��v`�9��k��O���clK�/����ǍN]�%0o=�`�W�W\�]���͸�B�z"�\���4�;⽀���x:�*��xbK�!@����O��I҅�x_��$������(�G��$b�0 ��'g�5ӗ �!M���`�!1���]�ozW�SM�k�����k��J'�	<I��yP��o�� �������Aꦵ�ҊrKKr+,��Qi��e�������)�	��Q���e�U���J���;����)|��#��/vo޷1t�؃�f��<�v�|�¦k�6�Is�[�k�d�I���8�0~)^o����z뫰ʲ�Vic�(j0��&�hOBT�{{�~˂(������a� 7�Qv$��2�����<x�d�L�	T�� Gzy�ˬ)i?�g��e�~+�=HVu�F���Na����W�g����sŸM�ĳ�|��\�o^�IaY� ��K"�O����m�\���m�~�/�H�V�����H�F!T�������;�G��#yBШ��75�嵻#�Lٍ(�Ώ�8n�A i{�J�c����/���.)pDF�� ��,M~m$S��~x�f���@aZ��b(*i��պ����yO���5|G�5�~g����,g�m��m��ϵ���i���&�x�O��3�"��Ӯ@��;��f��NyUuT��#�H�n]�C6C^�0���Z\�b"�T�[?�+_�=�� A9�� ���g,}�@u�1(P�DU���s���.oM�'"���K�ZF�A汣3Y�p�q���Y'O�ݝ��*K�H#�[��G
�	j!�eѕV��OIHg�]A'vvG�#� ���?Ŏ4J�1�3�=�h?ga'�.U�@�H7���:{s��lY��fIXY�]GfA�R^�^kr$��g��C�K��#����b�0�9�����|;YY��*(�б r��xz?~��2$Z��,�$L*?\��W	�[�h.u�q�n/F�0Ji��v������y�u�������`~��	�� ��P��Ţ��+�q�(¼�
üi��Jtf:X����e��A(���7ю��O����	����Y�t��T&���:��XFR��|�͍_2
�kl���y��'��=�R�j��-�ʴ+�)��W� �n�m(5�!�P�C�~�g��	8��G	��t�wl��D9���8��7�\��z�W�8hr���pG#T�DDz8:�s��/|! �n�M }҇tv����to�n�"8s�Nkl����_��\3|R�
��C 8��d���ug�%(Ȝ���&��lE�6-�6&6�&r[J��)kװ���q�OC3ү�<��G��㞍A~���p���~l
�
/ɿHih��g�o���ehictP�����F���"��:�Z>	��%���H��k+X�,������~����2D #
e����<�Y��b��E��N�]R��[�9޷H�	�#��G�����C�	���/-��M��c��k_���,K�`en$1=GT�3P�`]upd�rcO�^�Ԉ�bмtq��f*�+D	�7����>�5�0d�5����=ܩG�f\�~�	�e%���5��s�::�LO�!��ee�E�C�`Vhm�*lz񯘀N�a�&r������Sѳ}�in# �5�����\�zQ�|��﹨�E=�o�TU�|�Rr�ں'<�`�:���+���񆈈ދ���E���g�k������NQ4�O3Dvx�}�.� ���ׅ��{c З�6=)�I���bW3Q�!����7��?�Y�H����� �����'�3b1�q�
�k���|ї��3Z�
����G���>3�z� yW0�X���I��|�gA����Y�C����0���*RݟкVm�[�pj>)����~#�{a��b����@��"if�ZMzh�g�����5����)�t�	j�H[�.�-�u��3����*A��1u)zQ?�5�FX/gE��-�0g�X%Sq��A-t�
7��,^W��ǽ;��Y%j܍A kQ��yU���5�4��Z�Q�^�;�*�PF<�i��ZW�ɮ�mt�N��t|����]|�e���=b�5=�7��(|�Z���z�SF�Df��⢷����w���Sn��JǛ;�wCF�l����=T-r�qx�8zGS��f?�&(f��KI��Y���!��J��C_m/�`UE��]�8�u��"MƑ/��'kr
^��m�'����뚖����E&ڳfdK��\��%��KC�-AGT�+�S[��D�T���3�f�6Nϡ�޻J��Z;��[B� j�\���.W��n���hv�������?g����3_��N��m$#R�H� �)�}�g1�i@���xM8K6�K�O�~�kG}��"t�ĕ�p��[���R���#�,jMJ����ŗ2q�B����
�7��s�":�x�N"��/:g�D�P��$q1���q��9�]�*	O��{衵���ZJ*2��[YC�N�Ue+O��e]�BZ��TQ�tA����X@(�]N�租J�̉������5b����g�	�g6���<����z��Nb10��@`��ㄒ�s�Ju�x�|N���fD^]�k�C�4�i���7�>M�9��il�xU�� �Y�������X"Sf ����c�?m?�C.�޸u�{C9��"�pX�]����N�i��HgŋlH`�uP�<�cL�	}0�;�4£���r"ut"lګ�'��S���	�y�L��a��+ud..�٘C����k�.C�#��Xt[Q����^C��S�g���lΊc�:��?��!�� Ȓ�Q��x�_i����ht���q��$LA��� 2Fҥ�`^x��eƷ��J���H�$��k����H�0Q�)��ԭ�VP[���c[�_�W�f��;��2 
�͢� Jc/����RȪ6�q�:��(�G��·?t�褑ٸO}3G�N�N؅q�,��D=��]�qe�/�M3X�Q��6t>[������r�j�*�U&��0� ���!|�X��W4۞�u�9��)��md��I;Hj�'���&��:�à���>�/OF�y���t)_ J�*K[�KH��EL���*,^�b�}ČYO�ƤEE_����|�F��A`���^x�)�ɱJδL�pKE�)�!�S�D�4_g#p��Q5֐Ew2�/����>�Ȩ}O�OJ���䚔��^��2��H#P����z'M9K�w;Ǿ������/�9�����������7�E�&]�ͪ6�K]4PV�۩O>��3Zj�s�\�a�`�·��F�^��ir��g��O�6E�2��.A�o�zW0�q�yq-���8��fh�H(��I�)٠`Ty�F�k!��֔�'#"�&辶�邆����k�h�8�*+$@V�kC׍�5��=n8���CjRX�@��y��\ہ+��ݻ��=��2��� ���	H:�y���Q�!wwأ�f9$G���\�V��߉sD���!�f-�����j�"�<�ܘ�&4V�x���nE`c3#����l]EN}��0ޓ�@�W.N�eҬ�y`��	�P�().�B�m>M��E���5w�gd����{����qz��N3[�"s?��zzE�����z�X(��b�u�� p�G�~�}�-m��Lʮ�P�[U�^�\z�W�_}6)���=�>O���	sD�Ќu2�Z<CI$㌏r/���>p�K�`R0�,�����`�Ο�3/΋���0��l���Q>�-���^34�a�]y����h�87>��?�����tb�_��5�qyգ�ݥ|
F���<��e�1M�V�~��:,7�3�� ��*ί���>�=Z�,��6x'��϶?p�����g���:�C�q��c�kb��t�Cp�G��駑�����PʆASTo���[h�۝,⢸4����88뚦�}��<��~#�i���B̛i���
jI��\�
�����\qkwW5�*���l}�!��0�dw)������65���ad/qa�.fڤyH���`-)��W-D��P4�+ōm[�Ԏ���K�m��V3�l3���$����*c9Q�ưs�8gB-�{�}SX�b���R��oFl7�:%yi��2�	= �(���*Ī5��`�#�P8�rk-���N:-#��퇖މQ����ќ�d�Щ�hm�F�Z��?��y](����%���6����S�BK��l�Q�N���8���@e2ũZO���b�h��cAp�����<���_�}'�i�������G�%��S��R�/d�X�<aI��6�x��\�W�h��+�BE����ɱ̋�_*���W��/4e���O���R��M�g<8�N<�g��	[�}�6����3_[���ف@%j'�\�o�&���"��ftB�k��}^oD3ֵ4f�.T�h`���.����M�
iյ��dg��*���qu�Ѿ7�
��Z���ЍĬ4!���C��ߖ�8��I!a����0��pb�����=�e�q�	v9ڒ��[�z��?��vL��~|&��1%L�]�Y�����&6�ӑ��s1}��Z,��H�QZ0Y��M��i�j�N}�����sM.J��T��z8�K�G��U	�h���G��#N�ɍJ����+Ɗ��(����*�[l�A��(vu.|�'	P�G;�V֔��7�G��_J2o����晊c���7z�HQ��&��?<rϜ� M��& A6d�G����+�܏���&�~�7Ƭ�#�E_x��S%������g��kd��ݾ�_E� o�@oGs��3��xѷ�W���w��jV���U�HZ���.ዦ��0`Ӣ�:��_%��w��l������7��U=t&9��\�������Ð�Q�u>�v'�3�M�b�	([�C���בL�����nK�p1s1A�.��y����K#���"�V��=bj4EuQar���nV�Ŝm�7�"��2�E�L�7+�p�P�F��8<�iB$�6COj�k�W��F�x�������85�@��2V�&���}�B�˨�d~%��ܠx���9!3�����;�w����(CT��n�h�>w��`����_ےo���me�Y�(IǼX'a��	�+�T���y=�--w+��K���S�����p�4�iD%�(�ʷ��<7�q@�7���}�M�W������7���Q��V��#8a�rǕ�vM�-��N}BL~E��9������!��^������(|<f���X������C&N5��u�q�H<qp�ߵ��%���%���F^�Y\�;�p7���'a�W]��bwO�an7�A.���e�՘�>?��.=8�u�ҧBA�-̥s��y)4<P��&��co2��i��q>\]Z��8��o=�n���v��+�s?���jJ#C޳w�Dq��Ć�8���삷��C��S�I�Oaz�WY��Zc���*]ФL��� W�mq���#)L#�O�G7�1,��A�~->�{yo(�E��?�_�7�W�Ͻ�ۑg�����V�S��v���~��7)��~�<�I�d~x��<����t�'�&ȓ���}ھ����Na-W|���B�_���-��P�Rb�=�=���!�&1W U���Q��Cg��e�Lo��^�Q�L��H�ܘ�F�A��{?v2������ё���I(�{�2�N��>U�X�I��������KQ�7��Hۇ��v�HZ��.��{��%��1!H�j�ڦ	&�"Aj�}I�Y�:��P۸E?��*�W��?X��.�:����]"	�� ���%V��4fޏl��L0�(����}�@��
��у\���~%�w�ƃ����G�qHu7^ϑ�����kIjC V��;G��IŐ䵮��#M�(�K,SC6-��c�<� �eM�������ם7&���I5�V!~��:=W��f�z·�~��^o�"�~Ś5r�/l0���^��	��t��x�.v.E7'�԰X ����:��v3�˃�茹�9>�6l��\iO*�LG�����Vd��^��Yd'Q\V!�"�/�~v!�yv*�T�ó@�y�=}����k?�'�� =���v��X<_��7ª;��}C�{x����Dڢ|�����\�"d &3�H���@տ#j�Û�b���F�EB�kؘz���A�;��1O<F��t�I@�#����zi 62r��١�O�~ؙ3\v�J��~���ڣ��~ �uq����a���0KD�Ć]�X�˳,����9���"9&�z
K���!W��M�.'F���n�@PK���/���yv�hN�����O�箯��-7�a:�'&.�7�s��כ�(7�M<OZ�v����h�9�F�1�4�h�y���W�wAKڎzF8��B�0�N�u~!$���
�S�$��~VQo�$18Uҗ����1	 `e&�f˾�����u�:L�D���)�ޒOΩ��V�m'ٗ3���tb�LD��������Xsb��=�j��{8l�ͼ����坖��fN��S��
�&�gW�<��n8�!L���X�JAQ9���h��KJ�M�Q�7��^�̠$�LN:rE	bW�p�u� �e�C�?��� �m�>�Frъ���B4=�� u����1b�N%c���2Ԭ�)¶�����@$?�����b�h�~ ��F^:}�sG<p�(���PZHo�%�����˯�߄f�6qR��&`�k��n9	�\�~�<��"�{����7�n$�����ѡ��U�9K���k2#�ݍE�ҁ7T�vz�rI~!�����v�n�K��� ��C1���S�b`oҹ�j*4v��9,F���qr�?�8�/zP�R:M���)�� �oa3�{sI5$�*�5ŀǽ8�p~�)�+������/h#�B�%��)��0�ݧ�6Nh"\����o��/Z�gn��/��V5{a}������-�KM���q^�_�[�!�%��!�"���("V�uD��];X9\��#
���F����X�O$f�{A����"F9�%�P�5E�?XKe���v�8/�I[j�%#pŦ�	��M��U7q��D��g�@����ix-m����
��_7��Ngm�wcu�E�dc��*ᜌ�a�ǥ�vD}�X�,���G�M�/0�xs��_�����^�^$z7ҽdi�����W �z��=��˴���H�����4�5E���S���dR+<~a��H>�@~�ȕVUϦmӮo����OF����C2��Y���C�I��h�Ir� II��_y��y�U=I���4�����:A���i%��'�4$:����,����,3��cҲ�x��������Xg�ꧫ
����Y���*��k�.[KJmtl�Р�T ������
�����Q/e;�ر ^�
_X�
����P|e+�1�m�~�â�-2/�3J4��Y��4;�Ƙ���)��[%��^M�*x�٘mA��u���(G&)گ\�od�I����[��(��w�r�(�Q̦��L�Hͱ��t�����_y�8�i�����]�Y�7��6�+�,:�F��u^&�F��,S�͋,�5�p�P����BAN_ϑ��g.	߰-�8	 X��M�+�j����\xu���9����A��J�"�N�8}�:z�B��G�͹r2!���93_�>�q���,%T�҃�XZ�N���������8I3Jߌ�9�iry���$��M�-=��mq�)U�V��`$F<%��N���W���(�>�c!��1TО���Y0C�S2y��"�Fq҉�d��xk��-�0�Sy�48a�
=wRB����؅��"us�R��2<�P��m9����T�3�X�%�W?�y[0��(��[�/��[�yuL��N���)�L��S̅�uBFH ��@�D(���9������x~`��[C<�y&��# P�U$��5��F`:�js�>��P�(� ü�F!��/��\_A��/t���A<�.kN�TF����ʐvK��Dك]~ |��z�`�T|�{����6��6�+��\�Q�%x�1��߿P���J�qN�uQ��Z���F������/\��Z�B8�۝�d�3Z1fZN2+r]�43{$<���!�\�wc �P�G30���Wc}��1�ï23�*-�i��(��¹�|L[�v��"��"��6�I����@�J�6Ӎ���Tǻgg�����_4��,�%)�ޫ�F��p N[f���M�A98���k3署��H#.��.���@�B�� ��V��kֆo^(�<�K��r�}�8ɔ
�DZ�����v������#�����g��Jb��p"F8�e�����Kl���g܄�m��Iԅ	F>��&J�R�M�5i1����~�a�i`�";\��6���h���n�W$���i�cC�k&��j��r�W`���
�#�}hЂ����,=��<��:���d�Vڦ�=�-��!�x�6��*��p�b�˯ܚ���n[$��{�z��B�
��S����Q�j�o�2��\*�vMΦb۶�Q~�os���7Qޟ�(�ª�,��òJcs�&߳а(3��/�E"��kW��"b�7Vx�߸��g���}.�~���9��+O��~)kw�~��(��X��q����+�b ;���sX��׭���4�� /E��sC�)�����/���[u�=�H޳�p��",�|�FFas���4u-@�G�h�����=)@���v^�C���%�!i���T�K��	
B���Ik�{��%�E�&v�(Ti�~��� 	/��%������
eE�ݔDП !P�ֳ���$�QT2�!b1��}�B7!M�{�^&�Q�U�8���_;J�bo���� �����@Ǆ��%�[P�X�=ҳ�=!Z�Z,���!��I����(�9Y)�B�(���3��ZE]�r1�+;�l`�#z�p�ӓ�$�������ת�q�8���l��$y9�X��y�8��5��� <�0��p\�0�M�7�!EJ�KE����J�\�� ��8����لW+�l�ɀr����L�i�B������,��3���8�Zl���:?|!��F�x�^[6�u>H�T`A|��7�{��E�lD�
0����S��\5m��Z$��Q�v)Z��.�Vt4gր3�;"2����6R{1�@&�<.���9��l���e����K��f��2�c�����#�N�P\��[`8%/�]�s���l�-��2��@�rm����}���l=d�p�ՙ�.�
�Iql8�8���A����<��)h��yE���HW�!�k�!<}P^]��6&�*H0W����ܨ��	�G�<D�=ьj��NQ��'yLMT�0������:�U�b�����!D��`.t�	�u��]�C��l+�#S���� ~���xn��9�b�@�]q���f}�~�&/P�m�KZ[}�ؼJ?����?7i�_�kɛ�{鋁J�J��q}Wka���g+�[>/k-^�k	z���=p�^6� q�YxG�Z���#$�c�5s'��S���t�rI~)�	󑖇[ė�����i&_�>��7-�fO<d���{�lłb��h�˴�h���1�8�AO�9�բ&`0�`CxV>M1��:]���ne+���8�\lq
f�xm�r)}x�%�.���`��:@!ꐁR�~�&�|<y�v/�t�1-��݄]*p"#u$�4
��l]^�asɷ4����)1�c�nc�h ���,h��LE��^��"?�AE���W"/p�uCI��H��{鑯�r-]Ez��9 'h��y���둭��>�O��q��<S���P���Y9���X�����˭��ާ��j�ǲ�-x��ia~ʢ>� 	s+���i�AJ���]ǣ�o�G��2�#(E�O�Z�?�#��s�0܏2���ׅ���I��)��Y��D���I}�_�%�T�M"�K6 kPr��� ��n,	.@�}}�i<�������)g��B#S���hmT]��|k�����5�-��iR�_�����k#�t�g�����k{y)u�I����/F��ʵ��]�9O',"V5���v�	f^fCy�(�g�"� ,IQ>��j�J�g�W��u��Y}����|�0?�}��]R����3��iT6v�X�7��{52q��\Z��P����L�YP���p�+P_����@}:<)�.�W��LNj�T�����w7��H`���l�<'�5�#�[��\4VCS��g���l���S C+?4�N�>_$.��6T��!�cX��WI�Y�'j�t�%��G�]f@�ڗ�d��nyPl�J	e FN~���#�.k��őI�"E&�F��Z�����S�Y����RA(�������30U��J��B��J��1������(�Ij�H����[1 �$�+�rBt��]V~;ߣ� P�\7��"�>��oz�w>�Tɴ�>�r_��_fڵ͌|&����r��rP�:��2��y�θC�_����=����Z�B��KW�����{z��!�D�&���G���s&/Q%zl}]jFC�vJw�VR�~�_qh�l���(�W{Ӿ� �����>	�P��s<�*j�Fi�,1��0d^Q��9���^���x���A��u�Ķ <�i���
�f�`G�7)�!q״��K��P�,�!��:"o������ǥ��Ğ��w�y���P�|�`���.\6�t�S�G�3��n����ŏ��-"��4�N, w7�`�W,���������l����:�,�/�_z�\�\	�/�Mq�t�}�QI܈��D.*-��K�J�%�#��{ ��J��)� A�����Ŝ�"H��w+�KK�5@ ����h��簭0�������Ŭ��Q���]��f&��H�]����/d�/�w\h�Wy7�^�V�(�Ie:6?^�ϸ�JC��Ϙ��`S�!���҆R�κ�K'�� {���N���T�ʷ�ĉ[�����b�8 Y?M�Q9>�ܧ�Z̨F��j����aeM� �N=(�	!2�g�|f�9_%nt:�>ڼ��&�Od�-*��M���U��dl�j�Qv�u�1M���S�a�V�x!zn��ϩ�^���B�+���XG��HW�еA�fI�L��͟�z��v-��$1M���Zf
��up���a��U�M;��G�����jj�"�h��(�۰���9�������^�C�r8Ԡ(7��{�����&�⺎JG�|i�&m�U�M�7��Q�/�n	6c˧�gI�����M��}��\j$q���3��'O��UM���R��aPZ��?��C�H�ȹ�: ]�kC\�J��O�]�?,ѽ>���`�N.ﰅ���#��<\��+9E�$��-r�t�#��	Kd��ӄ?[X��m�n����ܘ�5����Cjrz��[ �F�j@B�� ��
5ܲ��Z��M��A��޳-�3���2���� ���k����W�F��Zs�x
��^��£N����#)�����m�D"�|�,�V.���9Q�5c8wnS����H��b�k1�zz4�Alj=ڠ�`�f�k�~��|�|{��t�ߦ�e*���������1�΍�cل�+h��
��0���H�y˶j�"��w�	4l��]��7���0��B:�o��h�*,�U�b
��#��xu�\1��Elj�}DH���6jW�K���K��xE5AN4=1؈Er�x���F咀�lN��T���׮�e�G:�㾩���]���Q2��0�6��RL�+��dE
B�r�V�^̜��"B���F�^�v�Iq���x"7��
�Ǖi���g��a�=EK��]Mu����F�ޯbd]$aъ���+P�/�nR&l(�6�ȨQ^�ώC8�Tm�<����k��bZ�w�fQ�Q�n59�����Obh%Ce�	�+ga���4�ޮ�Σ��$8��M�\���;�?��@t3���[(pG��z�_���/E�pK��V�����[�}�߱	���_�[�#�^���  5�G��J�=i9I��;@�Bom���?�h*�kK}{�N7�v�v���ӐJ=��0�P�5J��*�e�8.��*ǐ(�]��s��k�o6�]Fz,@�V�2,�����upW�V�1��e�m�JxVp�*ܾ�i�<���r*z	�ԑ��s�Y��R�8�R��2E�|�-M��jf^�"f�g�D�(l� ���=q-���Q����ӕY78-_Ԉy��W��eE�e���fƒ�O�>��C}l1un�Q������c��MU��4����Dz��t�R�x���'��Im��ب)Te�G#��2����2��xpD)X���H{N�T����x؆��+�{����g���HQr@�D��I��~"3�X�]h�O�̐�d&d]BR7o ĒT^���N(y�5Wd��|p!Z�8@�,�'�3X#���0�*=�HM���h��#���E�>��l�����T"�Kd� jG`(����R���W���2��y~U7����9`e�� �(�W�$҂���b�4qfà{�6vK���	/ĕR�Ws�s�|�����'(�Yr)����ߟ*XJen�����6�������t�')�]q�1���v(*yv@=�2o��G�v�Z��,�Dn�
���Y�Iy�<L�x�iaA��>���*�E,�j4��nO����xK!s���ti��D�Sã�E؎6����9Y���I�����=u�vw$��V7(�D=�Gڦ�Y����E��'��ˬ|ǳ�v�0F�;�����$ޢݲo#Ι�l���X�e�r-�5�v�����Z"���.����e��Ǿ���<i ���$��­��QY�4���x��bi���:tS���Z�ns�<�M�C���Jw��T����l���Ş5ų��.�W��m1�*Q9�
�{�J�_�4S��C�]��0�s��ּE���_E��6�v�^���\������ԊM�GW�[���0�&�C_�c�l�q�c LTE�b��V�b��E��5�,���_�?�º~����P���O�^�sq�KMC.����]���Ӥ7\V����$�L��Z�_=H�W����LѰ�6Ħ�
���s�-W�(O�W�jZ�.��I�����my��g{.��K2��(O���O���a���*Ƞ��'פ�\X�h�Ig �h�X �!7��IU���ϭ�UҀ5�W
 �C)H���Z_�I."�d"�6���/$T'� �^'�x+|���A��IZ�<[X\���l�	�-�R����Z�*F��Q����k�D��њܢ����1���CWoSS�3-V�����4�Gd��s��R�b��zr��2��9��E��!(����v����4������x�����5�: p����/_mJ'Z�Ç��C���2/C��??RܫC�/��h}]xP�`6�3*��R�C+l�� ���jiH�-#tB*��J��S�M(N��S��GNXՇ�����HB�`�	��O�������"�2:��3ݯI_" �OW[�-zm�*�G�s�������m���� �:#B��I������Y��Ͳ�I����v(�U�Ʉ��/�Zt��#B���JS;�+	\���bU�#;%k�Ka��ɸ<`�G.q��2�q�U���j��_Igh&{�{;/R����i�{Gy�i��&��a�7ʪD��)��H7Lڌ�_6*����&�#��O+�O9ʎ��<�A���BKh�+~��D��OE<�����O(��F������Jܜ|�:���J�3]A�m�l(�<c���2"�:7�QG}��,J7k�fC��P���In}� vp�(����x�M~�0�.��?٨ �|�j%�����Gx��X�x`fF��I�Ktc���ή�C�'�
,	�X�~鋬넽�ѹKz��d㥹~��QW�:�þ��<^�,����%�߷*��o����Ӥ�{䉰ے2�HN���%l�qh�qq�ҫ̥�]�?86씦�݃v$�'9W\�5C%�}0e@�Д=q=�s�U��y�*{]ķ������[I�q�`��q�)�{��)�&��xB�YRD��P/'���O�B�&�
������<hz�Ƶ �x�a��ׂC�{v�!(�S�I��*T�K�D�ԯo�
�b�pÙ�P\ċ�o%/)��
g��K��yB����V��Z�����Um�Kt�)��2������;/�_i�jW���D\�n�^=��m�i]ǒ�Pp�Z�V��:(ʮ6�i�<=z�S�=��a�▹Z��SL��	��L��j@Zڑĉ!�ſ�wa���.�ݒ�5��E�{DH]ؾyx<�^�/ç
�	;���:&�Zk|L�� �[,%dM���_=�p�H퀋#�hN��7��K'P�Cr	�g���T��T�I���!y�俞�!��奄b��h]���S�ҺDh-�Wٺc����R^�TJ���b|�=P(�WZp�u���I��n�Ӑ���T�N�Z���M��(~t�ɐ�̐i��N�	��"f����п�FL�/x�~+?Mʮ�� ���P�k9���Bu���@y���%cD�p�DE�� ���;n�ˎa�p�S��Y��̱��>9E	j���g�-"�"�؎}$>Neg;���Z5�8/2�����a���9�/2SxӤ������)��Z���"h��"�M17�(� ��1�<��=K<��hC��'Y��<�"��6u��>8���i�e'��np-��⠱`2BD��I����P�4�>8���+��" >"ͅ����E���l�����S+���:YS_	5�$�Uds���1K������u�����Y�%��>�=4Q�_
N�0�mV�N��F6�y���(S(�� ��_ͩE73f,#�HgA�7ԟvW��	;Y"�ev9ֺ���y�� �0�m�l���/O+��G���?�ӌk���>�v�@��*��A&���e��������+�w����?������Y@��qp�~t�Jc�hR���!�3��H��l(�B'��P�X�d(�?�0��(U&*�ѹ��BZ��4���-��z�A�̏,��QV��,,�mh���5��=t h��0�`���Ya=��E.m�u,V�!�ֲU�f� ��8?l����Z�.�>�~��D*㙈K���3Db'췣~B�{�7e%!��v�(���ʹ�ၘ��_j�6��)><
�t#���:����#*	s��EQ_،�N*h]Gٯh��-���\�ܩ�mG��L�N��>�{ò����U��<�|9U��*A7	Tmt���]���oh<�s=��� O�P��>�i�8��?I�f���o�ߎ�*ɷ>��y��0�}Ɂr�VyR_�&&�3�w�[-�eLPCЧB:p�ˁ#�o��i%D��T��%t4S(���?ꥸzKg�gd��!�1;�����+��| �{�������#вfp� �[��r"\$^�����7E�C��sFVǆ0I���o:ѫ�FH�[f�R�Qy����ԉ�"��P>�.�_DU���/�%��z��OX�D�u��<�O1북�3��͘^/��?y)xi�g+�L�`a'/�ա��p����U31��Ę��p�kc"�W���Q.����F��#u�/������y�ܹw��`�1fhN8v(���FZr�Sjy�bL1�5x�5�e�/�h��͚�uЗA�JI"A[.ȟ����Or��:Yk��P���}'�>VDh�{b�(��y�]���:`*u)4�ۿ���gZ��Чs�%x��E�" a�hZ���\i�E$h�DI�lRi�<h8��75�X[bk��y� �"&c�ǜ�y��u�r�~��e 9����/��6��CoN�eO�������3ǵe���%��]i�%#�����r�؁�����mDj�x�\y��ܙ��oTӢ������P����d�l<f��UE�io`g�\*J�o�&�J��<0&��r�&�X��.��[��i	Qvt�]%`}m��k�Zg�����\Wd��W��o2M�Uo�
S��1#�9�)D�eN=w���Rv_Z�Fr�\�+�k`�N��2����/��?Ы�o��s�d/�;f� �I_IӀY-�m{�o�ڊ&��/8����Z憺�~E�j���������`�>���%��9O@}���/��m&2�>�:�5�I!�D��I(�PR�J��`�y�6=?�	͵��V�i��bY���x��	j���OV���a��� I�4��S��o��&3>;�z�=�R}K�{*�ȭ��8r�?��z �ly�yg4����Wu�9[��ӂ�lL�i��v
8.�&?�w;v�F�j��J�v�q	'��>���_8�v�����1J�F�h�"@m[mC_P���6ِm%���ˤkE��\)���W�i�E__���6�cSs��5�8Rj�_ט>�8�"�-�����g���U�����6��"�������yYB�j����Qȍ%���&�I�Jw��z$3'��̖\����h���žQ=��O��6� 8K�!��R��fA�Dm�7i�a0��1�fJ�y;�����Ɯ:f���q�>�]`Eo@�?��k�Bt�3j���8X��5�-u��K�qo�u�w���.�ɿ%�u�E,@2��O�h�?����0b8lۿ	��JQBlX�A�X@��=Y.�F,�#��� n����E�Q ����/���k��l2���(�I�`x����}�7����R�!��گ,�m�j����	U�m}s�:�$)*��9K���[����C@+��x9GL�/oEr߆���i�Y~����
��Q�֯8m|�.2ټLc��黺�(��p�b�������q�.YfS�V��}4�.�ɣ�]=ڧ���S��l�j���=��g�h�=B�f�-�`�'-{� �LK��i�T����n��4z�WA7g��Tm���"q����o!��?�^�~$�˼ؓq}���2p�qkoAҺ�?%��Лޓ�1{6�P������[�����s��枦�J��#[�r���l+�:|���Hսη��F4�ZN&$�h#���a�^lm�_�l2:-p�o���'|�ڧ�Z`�w��{@�l��{S���(K��(�)[�e�4�Y6U�~d�Ę޷�o=�1�^W����\�K}ǐ��[ίJ\�p���n��������Sj�ɿ<}o,�����ܨ�f^|).�*��t��r`�o�����mo)�t���,g|�2V���4�uڒ�������C���I���>)Ai��1K�����	��h$�	�+�)�I�+�@)f��pU
?�Ϫ� Q�x�`,�A��h<�F}=�-�э $Y��a�9�����aRBh/�4aݖ^�cr������s���P��I3>�X��c5�1ŃD�T[�d4�R.?7�f�7D�ep\y�ļ:>���8ZGB9|�J�����W-+x(����!� ��>�hQ�V����xI����n�� ��;k�f��p��ɚ��O@LhAӀ�� �_ve�j�JA���BcF2�q�Z!�Ƚ����AEb�a�����g�!f4}�l�X�%���Ǭ ɤ���P��2�l�-�6HX%ՙH�<�㡨��瓨0묻<l̓����M�@f�R�+�B�.Jt��0]�~w.L���M���כ�-:=���w��+|7oY�ʉ����+�N-�''��'�F���ýGt����"-�EC]�p�L/��;�yք������E���#5����i�I&5"�8��[2�|w\��"ϸ�L~m����� !x���C����q%��������Պ	B���h�l*'չ�?ΐ���g�H�R�}��������ԥ]���G8�/���1B��u����.r^P��O ��L��@~\�8����c�&[�Mn����q\0Y ��2WW ���y����*�O.���#z*�&�}����5t����o���NN��SO�>R�S�ᬠ��_��ob�E�H�O������� v�ư�|>Db-��G���z��ͺ|��I�з��9�<��۫!��s
���"�0�=B2z툁fX�=�1i��Ս���&NC�F�jQ;҈F���r�Riʺ`�'b��;Į���u2be�K,y�X3#�-�N�s��-��TX�[�	]���w�:#���Pb���v�`�^<1�'Qo�.�Otoe�͙�U}�?��v�U�w-g,5�*/0=V�/�������%�\�������(rNս�M�f��d�S,��{��qҦˏQ*�ЇT����=�Twֲҁf�r�޻���@��ڧp��+)(�񢆯�r��xƒXR���Rۮ�/���c�U�(�W�YE�O^��vL�;*<�|@i����I?�m�x�x�9R$ Ui�:��EqQ��
j��� ~_�ך5niic}~/�m:�+�,ʞ���W��I|.�!�/����D�k RD���1��?w=�HM知v��R|�r�JД6O�ۺ�4�]1��!Ǆ��#��l` �n����5�g�\��,��r����k���������`���<4�A��x����D\�1n���x��%	�Ƚ`� ЏU��xP�v�!���N��>yAjq���5!�氊���u��l���쇌o��p�E�ʱ�p��<�z���=��s��V��^����UW5�*l~�,n#�!)4V%-��|���~u���O���FY��2�Tqr�``�"{k��Ƒi�]�p!?����	:�b��]雴�!ϳ�u�̗���T�� ��G���qQU���/;P-�]qҼ��1@/� i�40�a��[R�'ࣔr�A��s��|�Py�n�x�����"�WRj_1�q?�a�/17�uQ�q� ��f�Z��O���{@��ׂ��f�uM��d�^��7�� d�f��w?6� +�Yԧµ��l�F���9�E�*uܴ`�:=ۀP�����j�/�#m�����h����|�V����0�_ܶ��"�I�=Sj��-����Y��T�K�5������ݽl�&oIǯ�:t0���7�Īd�kE2�>���(� ��рUF	a�Kf�L!�mtpk44���*n䯹����h'���-|��f�<���wЖ*�Ѧ��������]7�i ��b�5��ʤ�B^��̔�%��]���TLvg����]#Y�!o�c�0���ڌEF�d66�
��&#w�*���B0սR������D�C�����h�e�O�ll���H��=��Ln�߅B���ʥ���5(缯�q=���Pa14�֪y3����ah��_���wL�!kҧ�R��ZL��y���h$��"�d=��' f/,�0��
.�YM
2����]x��)�J���(�mLmECp��d����(�G��̬@���j�4a?IA���_/��|�k1��K}��3���ւ�V���#��Bsq��L�
ly��-j��19:U�/�I�5x�I�M���(zA�����-�}�m���U��wt����aI䙞�&���O�?cb�D�a�KV����w_lD��vC|MO_�^���Tj�����nk�b�`�TN���ۯ]��ɏ������ƇQwJ�Bz�
��{U��*�ƋE' �e��>��V�1'�x�ي;�WGꆦ�:9w�ɭ��Og�Zε�B↭G_׊7Z޴<�^�<:��I�YG]M����c���8�D&#j؆��#�W�ם�3� ��o�K���C§vH���TMB�Vl�� \�*���z bG��9�`�.�Z���k�Z������."F���2���Cb�-�n�4g7��!
[EzRZ��vH�Ӌ���=t_���(�V�����D*+��^��x��;�\�~�}���U�@VD!<O�,oK'ӯQ��U���%&��T}�0mEg��ݛ󢲊��	{w��|&Cagn��r�1̗��=%��c:7��S􇗶c��<�Tq?�E��v���`�S�[��)s-o}!S�s�Ɋ!���Fz��:4S^��\w�u����U�d��OoNksf.>t�=YO���:�QM�V �#P���?�IB��V�xc�h� ����x9����^�yL�_��>�i�n��^E~A|,��dP�C�o����Sf�O��L��G��յe�N���	�Qk+���׃����"��*a�O�곏��U*F��#䶙n�e(=XC�jUA�8M���H�$ߵ.�����Ȏs���>Wݷ����곿;�[-j�P��)qNÒ��>����vb���}T�/)��)Y�k�^�-)���ADO
����(������D�L����{b����gm��\��3�F�eB���iᕹƪ>����Fӝ;�k���ɞ$�Ё�ٌ��]��b��F��\]��6�(3{miD6�)i�!���Xɔ��=f����T>�Tp�I����t���m&m����F�ا����xx���/��PJ$`�&@�]���m�p?�&�VEB�}r�%5nIF��֯���|i��&�lg�0u�o z6 6Q�-/���$���q?�[*^lA�`�����*Jփz$nL{J���Բr�~��/�j�������Q���$U��*�\�N����y?����U������ҥa`'���;lM��������5�W�k����*,)[!J/�]� ����ܴ�22��\s-� ��|5xcN4�a-fg� �^G��c��m6�L��L8H��|�\�*��(�a��Vu���_J������[���� �3��g��(P�)� �$��r�/:�/��%����:�_�Y�(Mb�i�����E��c4�9y^q��Y�����U�5̋w�W�|����BXE��W.�O�
�7x�d�Kz궹K� ���I���<�tP�#V-y���{<�����,�y�ZI�l[��^�$k�a������S�,ގ��V��U����bO�J���j�;�"�{ނ��)���@%�	�ϦXSdq�ZgG�*�$K���D���{y�ӝf��Bφ���RO�4�$j�j>ʱH|Cȧ-���yxg��*Gڭ"R)���j����X.{}�d�'�v&g5� ��E�9��_���gK�+=��,l|>�5s/ԃ��:� ��c�fe�w!-�d_hg2�DK$o���>�g{�8Ҟ��6��I���r���O@�囀���TbYǾh��\1��zb�_�ñ,��!�p�bsOboX��S��,�Br����N�+�%j�;W�ϖ�����{x�ϲsC�Y���_4����T�q'1�w���G�L���\ל���_/��\�h?$���q%hMC1�d�nl��U�J�zy�ۥ�['�e�&���=�<<�x��
ǂ�����J�����'�6D�n�|0�]�K�N5V;W�_b�z���!{e�z�.EVN�����b�RP��p�VHp"�K�E����*mpOI^��GX�IƬ��,ʘv����%iΌ�kmWV��nF��a���b��y X\���M�
.� �P{|��B��
�Z5]@��azh+������A���2��U��*}��O��fD�Q3��<
��V�8{�k	YѪ!�/�8�5N�s��qe<�������h&�x� ���k�#��&�H�����c�(u_ND{f-VG��A�`>@�6��e/iC�n7+�C,�gc�ƛ�x%�ZY)�ˍ��/M�5���[��̃��3\�kM�ppIc���p|ٹ'��o����͐/��%�:��v$�ֿ���P׀wt�� y/YN��W-�!	�A��Չa��P��ł��w���L��/�mZ	���H�w�]���U�Bn���� O�X�!!ޗ\��?Xy�Q�"�Z�ƱT���6�9H��!7���Tf�#wLc�g�U,�*��ob��u�kQ�J�V]����צ2����t���OYc�������E(=���7�c��+�wG�dlݲ�qir�3�h���J#�ޥL��7��7����T�������{��b�`�r��{�:��c��ѥG�v���{�d\4��b�ؿ:�(�(GT4"U���?(��ҳ�ƾÔgٰ|�^׷ݵ8��1���L��Ѥ���3�>:k��r����F���V�֔�f,Xp×sZDV�)�*_��@eΦܴRKښ�&ٜ���Ő>50��M]#P�� �-&�N�,��QŮf����Q����L���9vsH8�+����,���,ݰpNh�I�-<ג�m�/q�>F��nN�u���iK����A��(��_c��tl�\%	A��N��OHxC�A��%i���SD ˯- |�ݣ��
�!�굤����8���;e>=I��	V?/ �T��(˹�
��ȭEb<. Cڄ{C��!�ēkW i;�۶Y���S���v���lU��v=��;`0m(�M��&�I{*� #��t9)�����Vڌ��Z�iJ�m��ly�+�,��,]��!� ��.5�+0��4+Ns�,����y��~'2=�koW��q��擸����V[�L��V1�� 4=�!�"�{@"���)�z�[��0)�<��5��s�W�t�\� �c���^��o
�:Z�3�O�� I<��!�w�a_.8y����B)��q����5qt|�`��Ͱ�U0�B�}ŌA}ۜ�u\�Җ��W⡌L�(�"S�L&9T�뗬������<���c��qh�NU 5b�e�0Θ��!p�n}�E؅�[0{[�kT�� ���xKR�	���B� �$ZVrr��E��~�PsGf��@�}�W��9t�=���sU��_�a����!�0��W��S��񸋪�3�?^�zmn�`��W���eVל����`Mù>f߫����f4/P�r.�ģ�Ǖ�NV,p��rĻ�	� ���H�fx�'��k�4�Dک��Ž�0�+��S���BN�N�����s�[���|qF�ס����o��q(��+����{����-��w��LF�IvMT��&����}7�"n��b����_0ՒB��\,�e��4��qa�<��b��wWֺ�W��2V|D�P��G��2��FZ��:����N��9�.ɒ�M>�FCx:d�b�\F	�]��dt»���n��2B .t*�:�a�ϖ)�&W�c�
O�1h��F%W]}�ƞ� ��dJ\F��f��^�*RI��x�	8a�q{s�FK��{��政�����U�ZL`�%���`�y��O<�I��9�:`X��'~����Ig�� �5���ذ��ن<ww��^����ٜl�����ϕ9D�l�r����w6�Ev�D+$np]����~�)8�E)�̌i96��sR�D["C�X��3�7�ݞK-u�F��n ��W�6)TG�JB�96��^n�NY����ӌDp�|�SdZ����6�ӊ?U�TUb�R�9	-ۮmk�dQۃ�A d�(N�kR�O����W����@�J\����1�L
Dh$J�����e��O1�c��.�p��T��&�H;�&)O��Ư��A�v���=�PI� �Z��
���hwٳ�9�{w�	��iM4�o1����	��3�2G�4��tSL��͹�!5��q�+�1׈�Ԣ�����w��M� l#����0Z���C�񻔨���~�g��J�;Z0�e ��ܩ_��ZzU=D�rO,G�CI�W�Sw����dٵ&�^T��Ơ�Q���apۧD�LH$Ě��:R,��!����7��E��-��~必��bN�Z�; L��*�rjM���jy\i��Ï���zun!�^M��¦pt��oʉ(�C$���V���ṼR27����P�
���+8�g�0���$X�ߴW�O�A>I����G�r��s�2�62��NF���E�IX��J�_���g0��$D�>yp�/X\���O�<6"pT�0�!x�Fm(4������������k�;\f�<�H���9?�ު�˱sk#��A�g6j�<�AM[RVj�r���G����#H3���q}���zL���l|���^��E����:7�c8T2�u������$Y��QG�����y���h�nO؛������5���/�ҭ�<�Cmw�ĕU�3�whf��@�x����uA���V��. ��K�(j�7�����3�r��`�<�>}b걾PP�<�>��K�r���J�^�JXB�p~��V]���0�=���)�T����++��9�������_��O��t5	��f�г�=���ް*h\l�l�J03;��+Hv����_�%y��g�ğ Ѩ�613!��O�c�bgB���V~pbe�I�XR�;� �q]|����������u2#���4��3L�x�Q��Uh�"���q8��٭�Y���
�G�Ɓ|��S��|m�c$?SIT��k�$U�h(�xUm>x]q����΁�j30��-F߯�7����p��٩���G1S���p�R�cyC�7��0�����3��������ylg^�:�]K+���L�_O#u��{gJ���'��?-Y�)%��t?���D���*\!h��� �a�	�p�.��j��^^��'qԾ���蝴\Op'9D��}C����d*�؂�^𓻨5R�"T����{v�y���>��͞�RV�f���I}�F���.!�������X�$�O��|~RU��v���>�36TA��|���֤d�s����?p������}F���#�xsi|�n��gZ�0Z�1�d'
Ji��m{��a^)u��[�Ӌs�?�/�C�z��n�k|�+ԟ&u±���Z�
!8V&�v+L�
q���E'���4ĕ%�����/��Cf�;�h9Hp�D�c����}.&�3����BǨ�����O���Bg)JjGd��Z$��`�M�Hq.Y/�}Yd�Y��	�-m�#gl��:��*��3ºJ:)� QBŲ]����)5A�m�o,
�
=(�B����S�潣�x��3�뫡���PE_j����uiR��S�ʍ.7:�ڻ��{.��T#�+��UV��/�T,]iK�v��w�%���+B�i�P�6*�{}�Z�����QP|�C����SDr.���И�>m���
� ��������Χ4�9a���	i��+J)���<����&����m��m���T���1�p�{���V���#���Gb�W@v�.ty
P�(4\���I�
N�.^6$,����d���2��
wE��&6Y.DT~Lvi���<�!����K���P� =��X�72�ФL��
�2��3���z�o7�(&m�/ ʪxj�z��;�T�+
��Q>�np0L���4��6�"��ál7s�J�[�>�YbH��S��:s�s���;89����������H�+��렚3���DyE���e��y���ä@z��Ѡ/	@vzy���y�q�n�G��t�~�\rE�e�#9��*�c�'�n�#�هۥ�����"�\�1g���&$�R�F
-��J	%;��L8?$-F�r�1�"�AIU��P�nA�~Yrb�]-^N��܈��۠�R���p�6�ŵ��]�a����+~	M>�iG/����ᒍ<BNr�}xm�V�.�X�6Am�&5��o<"�b�!zx��s��`=킹[tMG(��N �J�	���L$QM��ŹMki�G�Q,�h��tU�F*�O��!Du�*3{ۦ���K�(�^8fr���:���o5ᕵ�:	:�@Y;iB��cnh�|\	���.��5yݍE��t̎���%=^H�"�Z�ee��H�D��������=U�d!2 t��up3����:�+��X|������Q�CѶ~;��t卩&"��]V�)���2�4���n�OP �>��RD�����+�O�ѐ���G��w��>���^B��F����ۥP�Rէ��6[�<[u���jt�Mvk�1����c+ P%;�35
�Rg 1#�耉=Odl8��,'���5���l�c�ڭ ܍���Ede������ض��(�U�3����0C�L�c���DӬ����o��it��kQ*ٌ'�b����C
�x�T*x����u��Ҭm �S�~��'$����1r���*!���ax����b�7)�e�4��j9鸉T���r�͉�ެ���ײ�H�gM@������m�>(Za0¹�jn���@u�Sl�K-M�{l�r���c��QgP�!�q��#ܼ֓�6��x�⛩�Y� d����{��qlg�_KI��&���OX�8��o���tPc�q�=�\r�y�qS��v��S5B	i:���^z�������A�;}��(�$q��
��h��,�O,g��lSJ^]=�u��8�E&�aw4X 0���(�9]F�YG�V�-�p��L,�O��P�!�����O�]ڟ3s�͊n)��|���ER�(_%�Z�,� �~�ܴ��Z�����%�M�ظ��k�x�������=_:#�B�H ��\aA�h���������ɦtR����iQ�*A��jJV('���w;h�H{��\ ��/c�6s��jt���0l�'���l�E(/o���(�Mv�=8�OpNC^?����_UN��fIءI>��%���:L�K�Kr����eW��Z���B�x������b�C��~^�}��n����ΰlX6�FY0}�4v�ÂU�eS��_r�Z��0%���F���;*�.��ul��EI��_�����`���)��`���~������d$c�����ehŜ�^6v�+C�0j�l}f)���@�ϻ�|L���'^�΄m0X"y�HŘ	�I�Ifvġ�ҕw$_����SbQP���ѕ ���A��b%k]��a�O���Ʌ���^2P�%�v�N�	�.,�}k��e����&#cί�Ddy�H(Թ] �l�k�[p�8�?�z�ę-����\�A�T�o ���,=8��0p�q�ӫ�}6y)<��n5���Ż#��{}��ա�y5�Q������.1 \%��M{���C1�YrΡL4�*�� �S`�ʇ�	��~�[��x��#/��w8w/ ��$l,>c�'5	�Z�_R�4�qj	'��!��}i��!Q�!�V�]��FYL�*%|�����)^ޖm�t�T�I�6xӇ�`�&)է]GW΄|���q���-��|ui�tiX�#��Z���Ha !�&a���"a0������2^]��&H�A��蔞�`:�z��n*�ձ���N҅2�d*(*�?kҙb(wc���r����ֿs땔�t)�$��(�xr�/�F�ڙ�v��s����Y)�(�jGB\.�M؞��|q���B�����c|3j64��e�����#��_��{�	1��	c�*�x�IY/1��0���	�j|��R����S&3a�Ly�|��{�_?�t���HkVבֿ��wly[`�+�H2l<�T�U��!ë	�/�W���JS���H�ʦ��?�u1����9�	���Cì�q�	Yl��E|��f}����@�A6#a��7՛�L��dkFh���~"���js��1�6���w�}�S�}/�D*��Z袘]r���Ӆ�(��σ����+C@�Gh\:�A/�?/�А� '������{�+m)۳���2���h�WAa!�b�I��t����*����%�
��G��G	�ǽȔݡ3l	F�E"�N���>���k �$�&�TϠX7����fpn��i�ߖ��V�h��4x�\9 &�b�t���jm"�d���"b@�<�Y��D���b�����$@���P�th���y�ߌ;�M&��+���J�� '̂'�����V�q��+�����^��j@��O�wV��3>mQ)�*>����h+ȭ���Cߜ�,+�����4m��0�3�brq�����h{7!�t�7�r�kZ�	\Ό ����悌 �k��g�Z��{N :>���o��aBؾb�E�jɔ #HtB�qt͡��T<[���Q����'@)tC�T�� �6�C��ZM#��.K�E�o���/3�����`��0%e_Mv�G�bdj�/W������L�i�*��V	��;O�I�j�7���"R�\Ox�-?�՘+QPkl����Or<%+6�<ێçi�	m ���.�K��Q"��o!������%�D�*%�-�A��*�O�:>v�F�'��SSi�t@z��4��Mk����*r�j,o����01f-���V����"2���j����֫�g�jHOp�H,�YC�蟴()��r��F�����3�py�v��ugl�ø���<C�:+�Yh�DÎ(���,}���p�q��g�@4ү��'��g~3�r8�\3{n���o�,L9�=vKɨ�j/߹P�@L����$y��a� `����1-c�v����M	x�е���?R�D�e#.�̋�h�X���� ��@�Sj��Xv`�������8cr1�%���oN����X?G+�A"��'����w�\m�"6?Ð�u;L�Ǖ�����w�4 5�Ji��;U��DGe�VE4D*G8��ûGU!]�d��>+r`2�m{K�},�9Q	�l�"�R���M<��v&`H�M/i���*Iуǡ@m]��\Th.�g�y���g�̏Zk � �Q`
v��I&�pZg��nE.�)�p�y���0�8��FCm�67�1��ނ��jGy���o�M�M���t8ܨ��tmS�H�<MA��!�&�\����a{<��6���A+�%�ƠY뢬��_�x{@���}����UK[3���Gw{����rk�a2�(�t����������`���������Al�Z�PV IVmGƾ��m!��õ���
�� ��Z�ö��b��1FW@���߮8fxD��\��أr	e5�x~W�髡����M /�)f\�����T?�	�@/��I7��͈ѯY�s�� �R��ݙ�	�Vf��(s�>�]��a6�6�X���-��U?�Nf���{�_�i��9�'����hs�`�D�c�+�"�
��\9�����k�:#�g+%���5~S#W7��b�����Ѻ2Y���9p�c��;�[�P/;Yq,b<�*��5qg������=��Vy.bY�f��,E��k眮R7�q�7���!]Bay��׼���%�X�0xlZ��/�Y���;�7�`�/���y�q��7�ɡh�6�^e,�"=���
����v�L�Q\�"���yn�&ō�q��1V�'��6�OFD}�ouP�R�Iw�)�;���D�t��ǀ��J��.�H b�N�>�nT�Q�n#��u?����������bሌ�XL����T�?��tLS���.��%Un�I�?.��G��Y�o8j@+��iuե�� �m!$<�����AY3l������#G���σo(���BZ��bE��w*��kl�E�7?��+*>K�w�oR?g)�3� ��;�,�jq�����@�]<�|aX���g'�����q�1�oOh�
����3؈d�J)*Lx�2q�n����P�
�!� �tv=ݞj�B��5�l��07�U1���1��M�PXyuD��	��O�aB�P5���9�Z�����!� <�T�",��� ҍ���"����7��ͤ�L�5O��l2�ﮘOh�^�+U�j'�,-�>G[�	q���7�Q H�9�d��}�0a<>N�Ĳ��ܡ�s�R1כ�=\Jf��=��3�?ߎc���IJ�\�I7IN���LgMR�D�"RSk���=1��IFZvmY�e��dgy����]tu���{�>��T�P>?�q���Փ���A�f�
��XLJ"vN%NZ Yk���[�����b�H�&:geIW,I�T)�u�"\�]l�2���.J���ւm���Y��N�?����>N�ۄ�$�ȫ/,����2Z|!CH!UT_gv�o�E5b~���}�MO�5���@����g� ����DR������b�5�r	�� WM�ϩe>�i
�͹^J�{�֝�y)����X׭!j�=�����b\z���]��t�x�Aw�(�a-J�6z����(�u��v�]�f����$1'�2� �Yn!j�7����{2����cjZ���>$�b�Kn�Yl���17;їY�K�����7x^��՝m�1DO+Dk�P�Sd'�U����49PՌ'����zz~�𼅋�N��w�E��C4w�I��9��=*O���89��{����5މ����#1b�jjK�&���JJ���~}=0�=���Ԕ�d��<���eU1h&hb/�u2��{ݮo��9�y�7)=���%Ə�D�f�4	�8e2>�%��Զ��������>Li·�?!��\š��*��w�D6��y�Fz��LL��F/c8Vxg�~��&�78cT�?��*�\��#�G���]�?i�>����Ejr�D�� mܚ8w K3T:w1�|���̅Q�]�3�y*�����:˯��}��E$�,�`E��S~�߮ds�N���a�7�����L�L-U���_�K�ʷ�,�l>�fءM�:�A:R�׈F橧+��x���E��OC��o��y+F���(��b�Y����F�J��p�g�9vJҼ�Jo������K���H�a�J]����52�CA��^}L�f�u&1���$�u°-f�HG��g)�%�M�u��_ p��!�v��1W��|,-k��z��WA�	�
����x�-TU�ڥb�[Zbk4b��\�����/�pi��.h&>@�pxjĉ)��x ,jP0�ajju,K�~uh)��ٞ����m�& �!�ך���ө_[T����p�WW���n�}�k����^��ִ'�>���Ba�Y�,t}��Pt�����E$$���a�0�V��nn����ۢm��q��|}3:��8,�t���Y�k����Suv���r-%hBv4l[J�Zq�B�V�ui9~6r߽<�<c���� H���@��2�$�r�����ê����_���b�Q��'�ָ�^�yT�,4;�#�}� 9��3ī���Ny��*�Q��y}�)ɷ{
�)k2��	Յ�$0�.�'H���f��k����'^�O{8�X���xNW\�C}C���5 W}���?�N'C4v����<CNM�j�ٙN%����P��!ƾ׃��1e%��ǿ�8J5U�$�M+��n�w@�lA�-���~�YwF$E"N�
�˘I�HT8X�s�x�c-kܢ���u�qXm8�	u��A�k��b���k^݋Q^uҾ�~<��(��=n�\���^X��ɘF9���LT��h�aur,�����1�Z�1i6:Ar�����M0S�n���0{�x�+$k��L�hB6{�x�p�D��%�o�����A�7s���{�8]1R]1Ya�ZV�5��<cH2��0�0k����[xj��J��_�	}������S���@�?�77�{�,߁&sD-tlt���.��Z<�@� �_Io`��T��w稗��Z<�J����Y �[���x�R�9C��%:9�)����t�G�S�-�4�sX�g&<���ʐKdn�`���S7j�U)e�Xb�Db�v1D�H�Gve��2*[�B+�c�HJ� ���{��#��5:���훀���M)1��齍9���p�jCf�k*�'���˜�/i]'�4�I~*�ra�1�,VX�PN�vE���BkOv�G�2���<�觬ֳ�ޖ���Bz����_Ɂ��g��Z�ٱ��Z͐��*ɞ�]������o�����	�hC����Ӽ�:S`���������2��"��b9�����-K���B]�k�ڒwu��P�}i�@X��0��dt��6"S%�a�:������I�<@�Q�MǷ�3�"�{� dљϧ7d�#���f���j~�����Xa_�p��H�2��C,Z��7+*�l��j-%7lD0d�u	͉���Q��w(����fx��oG��yJ&A�
��
�X���u���L)-�)+�4E��7Ԛ5��Z����'DZ�pgd�N�ƒT���֘_��%ej��k��^��vI�Pb�T�R�W�*_@�P�ۼ�JlL���Q��-�O���/�e %�Y�G���	�V���$�M:��I[�<]ɛM�h6y���~̮�*�Rmk%�:=�8�z�]X��Y6~W�@���C���C�(8T}���=C����@߁��mL%᠝��*߅gvVL.�{7�;�Jb����#��ʤ[��Gp����=f�V���#}���=}p�4�-r�O�B@���ut	���j�4��{��m��)@��PeX��H�X��B����9b�@!LT��+�xR�R7҃.�_���+/u�#`F]�K�v�HC�xd�DAB;>|DO�Iy��?%"9K�S�s�;���5�j�R���/���iz����J�A�dь�f�A���C����3-������L_�l��4<g[����;(Z��g9I�h����zt�Q��@���1�=?ۧ,��۷���D/3���e.N9Y6�����"zb��y�~v�*��sB����Dg��=��U�6M&�w�%qL	��b�i)I/����+,�b�>؉νЎ��\��-9�7^���C=gb���lc~V���Y�K��m ���ׂ X������
��
4GCT���!�n;���Fp�\}�o0�iJ��n�A��N�����
8������w���[��23"�|�<�Q�H��66n�4�x��˽�t��̈�����>�y�9<OlɈ\#{�F4"@�ʼ���+���������<�_c�XB��~2��g��oOv�o��m�Cnp(5�}�Ț�>jQ�6��Lp�/�x�߹���M���ܼ�.
��'���( m��w,�s}���bJ��6J]��L-zSf����\5������S�9���"52y�^CE����i})�'�Xؠ=��9u������zj��E]�C ����\�Y,kJCO	Џ�in�D��^�ZY˞Y}�1�L��̑K�8�Hm�M�	5M@Q5ZR�73�pUS�'h���^�f���%��T�`r��%˯(�nq�|�}`	砻�,�t�FF���чc�(�K?]�*%1�>��x����Ǡ��D\�z�o���:�J�lN?�o�#�nV^-�[��A�x�M"k��������h;z��E���?��uDC�+1v[[\Z��E�������p8
R��cd�C�ا[�/h�QՁ���mr$佳���E0�8t�\�B�$��lR�$��#R�sK2�]��cf(�6��
N��$��-	{�R�M�
I��*0"�ڥ0wҞ�0�("���R�Nϟ�5)|�q�=�0���"��K��:tZJs�E=�����G��ˢ����y����ػ����;���*�,����A�$f¿,G�6�X<�_��"�q�X��+y�Hb��->k�X`�A�y��+� �E�O�v,ᄲ� ���8H�z=�g1wӑJ�1e+�h?�Vw�4&~>�a���k�3�����sU7�Y3�����>z�@3V��J*��N���͛6S�p'=Z�o�&���G���أ��$�+�	�	k�Җ9ت���<��(cWMʍ���2����;��F�=2*f�)�J�u�x�59e�ӄ�$.��mo땼�����(?���t%A�E���4�4�؞����.���Ęd_ʥuOY��w�ER��n�h0�	���>"����`3&��&�`k�m�e�l)������PK��TU� ���  ���4���rP�O��w
��y�����@�*�Ոai^�*�MR���c��a��"���Ij܉��k�2Ǿ�;'N��6�ә�]��Kc�!��Ms �W�Q�2aȽ�7�y��O#�Ay�a�`a���';��+sf�G;P��t��N><bU+@|�G��M�j�� � 0$NE���x�@S��y�z�c�y�ɋ&T�v���#��±lY˴��*�&��@9.��S��D�U�������L��R�IZ���M�EC�е���%��d�b�5-"QP����;���,A6Ϯ��
MA��XmT�$L�����i��׾觤]k���Q��
LTh�®T��B�7�B�=�z����8����;�vˌ{���@�cC�)w�)�wǫ�s�"O����� ڏ�ļf���5�\����v	"�;J1Цh&���=js�&��B�ܖ�{�Kĺ�\)*��ZO{M�CKw��#R�Q�t��νh��	ܳ���m�}���e�xA����B�=#ƫ.��D�_���2�gE���OTg�n?�'�|�%T �n$	��һ��w7!�I;=tS�����g]��T��2�v�EV9J�y�����	�`̺�#�	���o��J��8��1�i*D���=%Z3�o��)�S�N��9��{!���V���xӱ��"��>���r�b��9<���bn��QwP���i{��+��&��M��k��.2���?n�g`�Rڀŧh̸��q����nWr�scl�
�j�k���=��t�{�(�!(#2�AB�H��0�䥽�)_�W���|��i\J*d�=X��㳰sp~��I�|Oy�s%�Xe ������R4�R�:;&`�����B ��*�Xa3A{R:Gm�q+���D��D�i[�۰�?������f�<�x��X��9ɼ\O�>_���4UU�C:Z�"Q����X+�@�"\A�����{�:�e�P���G�I�eD6����_�ا�V[a?�,�M��vK�+Kf�⬛�앍��]����u��eU��.��^�-G-Z�G�컨�4x�)Z���`��H�_E���V�I�.�N}l��]�oX��<Ŀ7E���u��b�2�M��˨�
-p-y���^������Q�r�@7]��g�`qģDl"����9G������H��?�md�#���Y*�a�>�����a��G��Eq?�Z9��BB�XD��8�Pu���³K�Ƚ����Ƨ��!��%!�<4��>\��$���������ۀU=�E�_���<�N���XpDB�)�>�o	lnWQ��ym�2y�\,��a�:eS:S��1e�\ջ"��GT�-�ӽ�^�˿��c��G�rZ�͜'���C���sOe���W�C�-U�_�A���B�R�0b�u���Ӕ�1��̸N/���>��]�v��
�,Jv�<���Hg5�ƶP�QO�پ�T,��"r�;2�k��$?�U��7����}U/�ŝ>:��{=<���L�<%�[��s�Љ�+s/7
�=M�k���6�Ѡ��-�0P�N�wئ�G}ص+��'����UW�Q�S���[68%M��� ��'��w�h,tD��41n�a�ߗ�А�]�1.���^G�G�{敠�"�+~{�ú_Ѹ�A�T�܋�0U�W�Y��I����|���S̶��d�`{b[��U���Phc�ی@�9sN�"�̝qjy 9>�%퐝'2/�Y7��j7r��?�/����z^�,��a�����w&i	�X9g�x"cb��q�b���M�8��[��F� Y��%
r� d�ӳ
�}����~�Fh�z��m98�*�	����@6�]X�KDr�]�7(_��<œ2}��/�E���w��Ȋ���l杸k'�SA�[e$���RX[}w�����Юw_pm9
�:�����E2~�7F|�g���|S���d���J��d���ؐ�E4h�� m/sϦ��itn�����iQ2����1<�&j�uiQ�Y����L��k�����qE���P���NH7\��Y��܎1��y�X��p]1�2��|��gQ�u�~����(	�ѩ�X��C#����i�C��pL���>͐A���T�u�t���GI�G��Q�>��������ľ5��4in{�|E��p���̂p���*���o7���kd?P0�x�_3��?c�=raW�L�U����J�M�(�������&R�*I���[�~�ٺϪ�]�;햫\���]��nA4��S8z�S��P�2(M&'�K<�fy����Y��wC�M��O�#��"*尘$�X�=���Δ;s2�����%L6WC.�p\ޜ��^Ju`�\G���$����#A�#[)k�Do��߼2A�*�z��9_B�H�����Ɔ��r���-��go9���OM�ah��L/�u$?O��2��!v�|�) }���۴a��?���p�i���p�e�I|�u-?T��v M]1�յ]����F��Kft2r�G�%v,u?D��������<�,2�D��A������H�W@>�؋���	�*��>��{!�V�T�>Q޽��s� �l!9꜒����(F;��LE�'V��<�:L��}�7M_P3jT�f/�1iJ��+J���')�����c��	w�r��Kn�sa�\p��^X/jɰ���BwS�T��!0��KV�	�9D�-�ڠ����RXeM�q�P�(H}����)�y�%q�c�hPmS4~���I锌�>;�T�G��F]�E2/��2������c���/�f�b�zrڦM%����=���MPJ6ˢT�t�˄汼J��sP�e<� ���_�((vL���s[ZRl���K��������T�TC8��V!���G�]�GD�| �'sb�ϖq��x��9��)װ����&��/(�6���N\�K�E�o�܌�<0�0�b��m��`��(��)o�,o}B�IǼ �M݅�9����n��y��3�@W��u��[X���p�i"�Bſ�Oɻ}�<˯�ifd��z:��l`�WN��ъ!�Q^�7!3؋'�㥞�/�L�qj.eK�y\˟p�zna.OWF��هIҊ�Z(G�8�Jl��(���w�F,��?D�=/#�	�#�}L��nx�n�+$����*�� ����	��3³��2��(/��q�U�sRb/�[�����Au�'Y��զx��O�ܞu���R��*�7�4�1��rι֠�g�yͅ+o�r�,��us�֍��Fy����jC�ݥ����g��*���J��G�t�>�Q����T�0�v�U�A_���zT����o\�ݍ��g�ׅV�����D�2�֍�3�h�.1����BT"$ל���C`3����ihFe ��1��"*�gD1-z�%�o���U���5.�'� �޴,�(���?���;b/?�Z�Ҳ����=�m���<V�P�]�J�G�jL=����ez]�b��:$�!�$ ���e���^f�Dӊ99Y�1GiL��us$�Jor^l�����g�K�)�wa�N�E��0�c �-�tF��b�40U]3���oF�ƢҖrЛuz�������s���
3OF���{��~5�a�sQ:NV0��1q�p-twytG�qW"m�`Z�f*��@�Yw�+μ?3�o����r�?F/�Lz�}��6?���;>j*�V�������z�!N',���m˶��.�
��O(#�OO��Z�c�
t�[�`�ϳvyiy�M�����6���!���ߵ�6!�NR*[��S:B����3T���E���?�����2 T
g�DӓV#}����M� �h>����^��B3`��������m	\��"D�J��Pjy4�R�6i�jf=�:�Q�Yj�H��#Ȅ�BY�"L<bN{m��aA'-�$�8�L�[pxi#���[�x�������ŵ۳- ��vI�VSa���H7��Łaa�n
���.�`Z֪��J{����K�+���(���)�l�F`��m%�V�Y%�z.�����V!y�����k\�3٪�}�F9�>��
�JO�˧�F&L�3��	��(���39	��b`'AQ$����X������Gw���5z�_J��Hk��@�4��ɨ��	q�e��%��yO�\]����,}yL�����U���)���@cc�Sl%�[����GY�������~4�솎�8>%|cm��-}#�H&͌���vc��~5�y��{��Ҋ[�3(�K������v	kAw�=�����t�+��p�����mK^/'���h���M�G>(!ő� ۸�/��V}_�[,q������L9Mj=�������=O�,2�� ��o�=׸2��I�)+�O�\.*!�dq"ԫJl���ɉ��DO�����T@��t�S������-���D�Ĉp!]W�F��h�e�k�<�zU��D�v}ܧ�N!��^M�0,�ɮ��@�p�9�p,H�#�� �b'Q��յ�o�g����4,D_�@|�b�)�UjE�*Sv���&;�Њ�8Z2m�h*��������A⯢SM�ܦJ�~9_��(�0�v�{������6�+����vN|�_�ʂ��Z�L�f�w{���s<��'�}v3/,����.U�G ���r���4���;�����1'��b��#�h���\�h*�9�p頬,�+970�HؐƎh8\H��OP:�`[�L��R�u%?�ǡ�ϩO����.��=¡6a7��K�Ũ<*�?��%k]��@�b^��?uM�������?�i|�%�Ty��@�d��Z�:ol1��#���{tO6i��˖s���6h��x.��+��5��+�U	࿍�ص��Ѣ�X��@���Gw�Gd8�P�2�>���J�UI���{�)���GΓ@�{'8t��XЎ�����q(#�TR�M9E�s�	�7j��Q	�z�֎�y)����Ӓ��X��n�� �4��ܸ�K��ϖv�b����)c0�$U�%���F�`�zL{@�����[Ů�/0[hz����P��aq�ٖ�����r�Yl, ���i܇JJT�s�6GtaC�_Pa��3����F,�����
��더K�L�C��a�"�	�k��b���-���e\M���5���[�i���Ŋ�D�S}~ڛ��O���K�<:?WI��w�]lI� N+�_��m��;�</^Jn&�3K?����ҡ��F��[��s���*ܤ������$^�˲��<e0�4����M!#
�P��Z|�W΀_f�Z��I�Ԋ�ۦd���[h�	��ޔ�Xh��Ȇ���[͵.�߻\�+lsDǁ��fK Af2��2��,��읆��+�`��;&��7��!��c��9a'��/���l7I����ң�E�J"�� �N՛�Nӝ.�s@���RX��s;�ڃ�� ����)��I��'�OɄrE�����+1�{˭J���S�|0n"�z��M�v-5j5۰�T�xv��
ߵ��H~�� ��KќB#����r���D�o�8t�(� ����Z�NQ65l����nx�!6�F�Q ���&�����I%E��I���
�^n(k����ؒ�
N��T:��;,�n��@�S9�}��{�|͂\�:����j�)f�(�h=�Pj�<�nxYs��Qr��E6��g��4T�u
vU�/�3�ivy������ן��5a/����΂k{����]^T!���3�����^� S�''N�է��&��É^��X_;RcR!���@�V�G�l,`���*��н��n��~�nR�ú���zm��G	�EV_�����2���R����-b�%9s�]����QZ2�:�Xc�4��W����Z,�8�z���1>8]M/������
(r"����=u$b�w�j�Em��0n��:�E&��MGm�x�7�~��Ѱ2��f���ǎԖ/1� `���?�?��R,�o��L�^o�䙙�Y�,w����ތTa��7�Y�4�߁��K�q�y�J��Q!�aQ:X�n��u^1�M�n�j�	�}�,�l�o����&eBbLB2MG�*0pq-�vK'!�������)��i���[	�ސ/�5�Z�C/�p��o\��<qV��-����7ك>��!��?؃�u7	�&�_,/t���,Q�&��y�?T��<�J�����E7O�#Cؗ4�7QaV2�QD���|_�a�̕"�^W���$�S�L����(I��D~l�|����~ӽ�v2.�#ع���,,T�'u�N�0��Aa�#lGz��;�=sΆ!��������F���R-�9��B,���:5 �����Gqc�tև�l���}0d��*x�"aB�b�$p'�u����?j)��[G)|<k�}iE���@���(�2%(J+;op2X�|I������l<I�7:�ܰ1�^|e��Z�;�!��mu�g��e��`�h^�~��=��>]����S!�;�#�\�ͱo�˙~�Ӂ�A�"w�>�5]�}��g�`��'P�s�,0���:|�>��4��[�K�]���=
��eu�	@h7��ɹ��Qy�Α����̷�F�2�Kb��0G'��r6�u!!1	���둗NR%inHH��x��R�pE�Td�����h���Dh�6\����+:c�Qٿ��"eU#�	��Ev`��x���?���2/� v
⋪:R�M��ꖴ��)k�x�� ����B�j��G��.F$��=H��D�i�&��sU��2{�.+�_Nfx��֒xؿ�Mǟ�̰=c�J�sq�"N|s�|�S��KSs�k�J���HJIh?�H�uH�;����37��T1�8Z���m#0���ի�"�/�rV�_�͜�4�˅�Ց������vu��;ʪ��q>"�Ȥ���9�	2̑�{~~gN\Wz�\�*t��8*��H�u���qS��s���(hv��bV{c�@q���E}�h�5Y�[g����֯ �?�f�������`��fM�'O�WR���v�\�ۏ�5=7�iЮ���[|�O���b�����7_ zwXRB�}��G��^�\��n�%�O� �i���	٬�?�/m���j;L�^$qi�YJr3�2z.q�X5���8�7���&���9t7�0�9J:xNN��O
�T,�*ݰ�X�B�=#�1��?������ϊ�1bxx/��L�Ol��B��n_�~����T��t���{����I�3�J�548���0+��EЉ��l��y�
$o+�3�
���J�eP�d�ا9~-57�aC�M���:Z�ƹ0*�7�r47�������v���<��L��X滮S��
th�^4,��V.�����j��ce�	�A���n�Y�x`��<v����M;�r�xJwtZ ���b��^��\_9��JM. ����0dõP$���ך�� ��U��74T��w�C��z�mZ��&J�2U��	<̎��<���6�9�P0z7��+�Se�k�:�g��fU�����MG@΢��+�ޱzG�E�Uݳ3�����J�Ro�i���V~j%{���䵢Ť�TA#}"�f����8�T�P�_&_&1�3�D�J;�8�������.z���]�G�h�'|�h�v2�2>3�=YY��QC@�\��1�72A�+�چC���B�[ӎ�e0��n���_�"���e'Wb�T�R*��2��3N$����)�IQo�;QJa	��V��h�<:�����i�3q߯����:�����ٯ��w��
�U��S8WJK�\%�"��ܮ:$.u���i�_�W:򨞰�r�7��'�(�y�d���A���(��.�2ï������=F�O���c�g"k��������=����<�8��H6��;�
��-�KT2�݆8�c�,A���|����>�[�[Rz�)�Ry�p����b�f_~c�2�s�F��N��@d�w�yS)�]���7����^��Su�n���Eh��!�oߣ�zA"��7�N[�z��]����S�̀�w�-ۆ��֥�f���3����37�����$�D�>@(|��I��q�̟W��9��WX�f�t������kR�'Q�@�WD��|��$	�f��y)��l7�24$gB�p+��i9ZdO��枼-�+�{���[���[�NjO�E�,Xߢy"{l��8����, �m����O��|e�~���"HۍKx�����k����B3VUk�ӳ�9���
����C����jW��+�k���Sk�p�� ��;⟒����b�x��'��C��c]l^�>&�@l��V��2���ن��H `W���=bUv�V���X�j�{�����?G��)<�����`�6��mY��d#XCc_�|�?���U��8��E.fp�p�gf��G((V���5���������^�i^�޽WH�^��hE�,v5�f��6�lU��Z�kL%�5���?q<fױ�a��ߝ�^��^a&m\?�@ �]mx�����G+"5C�GFم��� ��
&�6ő�Uظ0]���0�r7������d6�QG�^d����<�M��/=҇���
!�
�l)��5�A���
7�p��� �i��XC3eE�eSZ�(u]h8q_'^��X��.R�4!��d�����J ]��s{����]��=GlU&��=�'EhE]�kF�5Cv9ƎfRI���1c'OѨ ����S�}���@q����$$��E?��6�����dL�9;!� �ޓU ����)
#"	ڊ��6x�����������N����ҽ?7$d ����pH�S�Y���z�����y*,������ӺtO��j9�Rj@�筟�V�z�
M�dMU��p��0�h�F��T�ǉ&`kj����8GW��"P��wI��Q���s����=�4s�x��4���3�o��#��W�}����>=�0T�|q"VR$��d��Ch�U9�{o~�'�<�Ֆ�x�.ك:���ۻP!.%1X�]5Ǆ��m�o�ү������+����H�=6��)�Xc������Vѣ
û� ��)؆K�T�ôl��^8���G#�����Лù�d�o�E�.+fz��N��1Ls�,���6G3��mأT�-����P�UF�R�GC	�	����G�r�z��ק��h@w��ijC�<$g�����k'G��UE�} o��sz�G�)k���($Z��h�-�O,]�&�h�C��� `n�. ���WH�FLI{ }%����yMN�#��!�+�z�O�p���4�r�wQ�ƒ��>涡�BA�eCF�Ppѧ�q�rb�R?_���-�%YfY�4�o�'��޾�Tk�X��t������B�=���,!�Bwf3-�ڏ�cN��̰8W84��&OI�16mU挣�7\��s��l8!�ҧw6�*G`<q�,�ۼ���V�6�Yݖ�$A��6(q�������0�����cB��d����ʱr���  *H�Y^��r�0������_�sbW������t�>/��mDw���!��2��HH+bwB6g���DGf1�A-��9�1ؤ������z�u r����pRΐ}���<�[�V��t�sK��/�Y7V���c��u���j�
���0-�3�H�]��=��Te0�H�Q�
U]�� K�t�q�W��-�8�>�;$xֿ�ROO�г�8np���Ul����{��B�w�����4V�~�F����\D��jсto �/�F8�]��1;��q	��=s\�}�\�l,7��~��������W�\��T�Kc	u����;9��h�5M��^t�U�d^5������c��;	[��u��Mx�"���]]�Z�8�+0 �%Ĕ���LѺ����c�A/n�z���>QO�ET����
BǊ^�v:2\W��L���Ť'�Y���x�
�>�:���%����n� �P�x���4�.*��^���NI�|�p��݇���Z\��0���W�T�h���͚����*G��p���1�ɸ�1]����RM��@�Ҿe���QGZ��*��OܞY$�K���r���\#?2O K{�Z7��|�'� �;=�&鯝=������fH�/�(tb�b����иy3�P����'�<s����]�5U�hr�Ny�=R^|�9�eGAE�ٟ�z�E�R�%����x�z���o�LFy߅��%,��݆Q��o���S �"���	r� �u��z>j� �(��G���^G��DdƆU��#}z1\�ۇ"�8��J���#��ҫ���7��-��jn�q����s���`OK�m"®"�On�� ��6G|�|��uYH�]���]�1UMQ�y���b<�/��Kq�Z%#N���8if�e�G�y��3���j�$���n�t�l�j=�e�H��Ŷ����qs���}�:��q�wh�8���M�� ����1#Ua�-�F�h��CY�{e�RE�	�׵��#�{��K!r�eB�]ٔ��~����@���iW��P�E!���'%����}w�}%ɾ��C���qٳ�����_��s\I�<�y�|pZd7�lw�`�G`^٣�?2��d�-��1s�>��C�]�F����U����i�8[�GXp�,6�M���N|_���qRWO��yw�`n��o���g�ྭ*���"	�\��o�DC�!K\����[+��Rq�fQ����-�!�%�����q�m��P욒QںZcc(m �&�����|��z}�'=��0W=����EH:��^0�|LF�4�>�"�MƄ6H��;�(v���UyrR�0"��f�eH��H3zY��Α�����^�6���e[�`�lJ9[��d�2x�t*��(��.j�*�\�`!��7�nt�T�KS֜��}��#h����lp�w���w2@_������g���2~B�=���b�@,��P��/�2b�?�ğ�(8[\O�+�#l7�~)���UfR��bD��_e19{��2��{��SzKBU�gE�o�5���OE�u\���/��pP�.�zM|�}XtA2��Μ�n��Ʈ�I�11�6N���g����i7�}F{ۋ/�c� gz��Q�aC�S�}�%B�ٚ���o��@�4��0���-p�v�_eP��?�8�7�<4��h��PL)?o���J��7�U�깧�8����tvWsl<�aQ�i��9x�K�������y0����s�����_r���.�����H�:��B	�U����k:�:_����>�l�zX�oh��\*��ℿ�L�����S���F�&����Fʼ^:µ��ɷ0F�l{�2�^ۓ��/��ޥĐI!��VBRc�r�I�r˭����^��< 2�C�+K8�V���\N$M�f�j��).�1�l�ma�ִn�����k�|0g�+D����V;�l�Lt%�@A�-+ݔŚD�e�LRC�S��q~q��DY�����J�`��T�FA!*��\<���������1�-�B,�l����n�g���c�x��2���HG;(���u
X���P�2��?BA����Ro�C��ų{F���,,Z|T����x���},1�O��+L�T3S{nX�	��7Hp��Y�IO��Woq� GkP�j�&��ޗ`2j'N�Y\��-�7mmԅ7�
ϫ�=!�J�p˳�P2�\ʺ(�5�eb\Z4Dl�<$
Νu�~^Ty���P_N�n>�ghtϢm�!��6�g�R���#_jl3���x��#���_�1-ƻ,9;aM�)�����z�s��~�)�F�_t���X�~ɰPP�iN��?m2��@%��`\W��ٹ�� =P�D�����L�,�b-�?<w C�1	QR��}����}Z�9�E��P�7���y���#޷���=�Z��h���e��-Hk��i�0��LAo�f�T�����Wl(��1��H J-�!�\��i{��5��~g�� ZxҸ�B�qh2{ūt>����Ҥ.dj~�4���x9�e*|yoF����%�%��-����m��^,9�A��O��/�3�ٛ�O�%���qvssTbpm�5L<�g��z��L&bU$�W�A[�0�� ��� *E�6�n�xY�)ԧ�%2�2�4���.��,�H�>��aC}+N�©��X�oʊ$��G����"����x��Rl�]QP��Eu��fҴ�؀e����E3��cp��yJڗ%Y�5�ǭ:TgB�_���L����$L�'
dr�+���<1V�Q-��D����+x�~��W��T��?�`��A�K�a���͹�i��8ݗ���v�om���K
cͳr��	��Z��+�GRu�J�V�����;��v��?���>U�k)B�A���9�e[+��Ѯ��Hv�*���1 ���x-V�J"�쨂ˆ��)	
"Q�s��m�Ao�C�J�4x�j�Q�7���鳻������Z�3�e�n71Ո"��x�Ztb�����IJ������^���W��%��=��&���^>��$��FQ�F�+�]a�����!0I�����s�{�� � s��4I�yl,/;vFJә�O6�_�b�'F�qa�Ƚ��YF�츋D���
���dۄ�%�R�-2��֏��8�KN�5�~6�iDG�J =�놙*��|�!,;����DUG98��	��^���BC���ԁ��4XAY*�?���u���#=N0_)�/I����:�z�r��Ú_����3,�W%uV��z��7�WS�����`�d��4��I���?�z�A	t��`,_�U%F�ۿ?eP�$zi#J	�?�3�0�1M7�v�Z<��/���ˢ��[<�Jb�B��y��(��������FJ"�҅RQ+�ñ}����Ǣ�Ըe��u�C�.�8���P��V��q�����m11D'����>�%j���4�mˈ��z8`�G���c��!�[֮��YZ]�#��˶��1�[�O��nt�Y���j�|Q
�	@n�т�0��SBM]��|~UKN�v�k��v��%@`��"�~jgX��
U�l��l$�:��w?�	oM�ۛ��������
����A�}�����Ruw�X�P��>��%W[2�ڮ��T���T5��j��?�r"�-�NVn��[���?Y�O�/u,g��ظ�;��`$*���AR���ơ7%o�m�(��D���|���?|'��IS�W��,�0����u)ݙA��r@Ѯ��� =3����1hS�q��������c����T.���~�"����̯V6�I_��~� c|���9�ubW�p�K�m_4m��ǽ�4z��[ׄcC �y*�:��&���,!�YA�ȽR2i&��#�ֺ��<�Ex�D�r��6�]@ౙx���f���1VX��><��~g=��6,`6iS=�`��6Яq%�tK�U=��D ?�O%$�ѳ�@��.I��A��]U��.�q�v�s���%��,c��_S�`�cd�m>"�$^��$��˪e0��S�C�j`8� �q2�!���Y�X���~?��%{m�����Έ&RYHX`4vA��lLO�up�����0S�K:�3��+�����W�P����/�{�`���E"r��y�l��8����M�6���g�I�2#���i��`du��#�����Ƴ�,53�XG0�<}��p�w�\.-Zң�?������[Ꮟ~K:��΁��5&m6�7�t�s�-y{�J6=�P�~�$n�TP�>t�����f���ʷ�(vg�+�a���K�^�&�����5��C��j�[OG�]��D13Ti��������w��r�N��|d�[�F�<w��G��~�T`����38�ٷ���G&E�|�`oP�d��m�j�W�P�e6G�׳Qf�	�4q���?Q�#��7�JX(��͔�ڗ9��y榌�5X�Z�u��Ľ:�X��v�bS�V���k��-��u�R�Q���Dבݜ:�O@�l,�����Q���9~�Ͳo���
f�|��HQ�R�#r�m?p���_�y�3#-��?�k�H<���
�^�E��/G:�B3Q�������E��p����S�U�N�ް^�����$o5�+���_)��O�?N~�R��'w��`pN��b�X���o'��jK>0�vhZʵ��ٝ:�{ϋz̈��T�S::p�ԓ�,��(7)��[�}����퐌�o���do��no����)��(e�<t5]�^h�"�ym���K֖X=����FDh�2�>��#�wg��u���E�	m@��y2^X� �o'@����2�0����R�N��c��1� �W��0L�����5���
�Õ>��h���� {7v!T�+^��	i� �h<	��P2Y�:P�+�;�;�]DՃ�v��0ԍ�!�!{_�K�pU�vW�g�7�0A1���� ������ɣ��㩡d����Tۀ?�>Ȭ.�V�V�NG�X#�IQ������v��D����,�j���Ű�?���"��Ee'�G�B����0��Z|��[�UI�>��MP��s���]�J3�/�?K> ����}�C{���7��[բa����k9�RK�ɖ��蘕�p�L��ip�юABY�H���S$��A2=��P3�Cc����8%������Bkd�8��f���-;n�$��Vׁ֬qEzت|+��G�%��[�7����B�#�d�y6�,;��������`��/���2Q�s.i����\t��\[�1�A
�́cߗ�L����7)���c���>�Qܢ� X?����������4�[�=s 95�*����������pςq%�%��n��j��Ƕ�!�SS;X1���<p����5��������އ�	F����`�?(�������"�p���ֺi��L���$��U��c��z� \����M�P�'`Cn��Y
К=%��<�Bٳ�Ъ�J0 7N<ѡqf�XOج�Ҁa�����?�}�ڜw=]3-`E�qۜ��	���9,�z��1��в��9l;7�W]AJ��t�AK2=�#Ft'��"�@�hJi�5�`Y2h'�i�Ӆ���D6ۺ�*�8BF9s��S5�XQ�L���+d��J��Lگ'NT��)>Z�H�|�8��*HD�)�>U��`��c�7p�]��ߩ˅s���(Z���`m���م=��N�8z�����ې<Ԏ�&��_'� ���{>m躮����j��y�"�2�DS����U`���$V��ȯ](Y�zP�%a D�q��/XB\�4���{r �����<Rm�c<~.5�u`�������p��;)7��7P�E�[f�zj�/$����_Q�@]eL�#W}��=An+sl���}ȉ��ѹ�Ž���~�����!LZ�ӨN���2�C�
���U϶C�"k��P��h�x#�{ch4�j���Ƽ�S������i��]Z,��材�����S=�aH?�Đ��NR���t��,���fv��G҂O����\��gi)5Q4*��I����IW����~��Ʃ>�9�� �S����Ir~��֮;4��!��Xk$��_��蘵G�1�+1�H��1��"2��� (�+jP��j�,���'��t:�7�� \�U��1*O��j*b��ݻ�m����jM�/+E�N�B{����ɳ���|�!Z!�gCzn�UTT,1~m}���j�Q:�jF�?�.�X���My,��y�
Lb�D���9,8�(ⳊEn��F91:k�U[�ۈ��8�!9"oLVR�ƕ��"�&�����M�P¸�?�O.`}� �LM�+�OCv��A�b�����`��ѫ�$H���o��j�ϙ���$�\ɍI!
MeX���u��"f��
��"�I���KG"��<��/�'6�2ʔ��o���ͮ��!Z�)')�G�Y7��ןj�>Yنςz`�+m��2�!��jX��]m��� ;\������1c�Ӓ��(�����'��ZU�-w���$���X-��!U�:vM��Se�Ɓ�A$l)_�uGI�\��^3��\��gm	[��Ӧz�l��>0љ!-D��C7�Lm���Bw�1��K	R7���G8TO��)z�p�}FI���4��9�5�Xq���� �ඦ�xRa�v.1�S��>���@d��aՈ@>�;30�׊$���[>q�X���v��4�\�x�����1��BV�I�7O��|
{^J/�K��$yi!27�|t<�VI�V�+��9�T��֩��ϑB����0��qe��=��SJ�U� �o�+v��d������&�m[W�
g�p�HI��&ڀ��F��
6f>��M<Qɚ������d�B�؇�:|�(�ƻ�4�xE��d���zY���j1��jY�1g�԰�k�fﮚ��&�C�r1����%��{�+=ف�������Z�ФņjJ��y�[��B���w�Ml|٪�0�K������+��N��ʇi%��=6q~S������6�������ޡ�=/P �,}<aw<qw�S�B���x���+*��ִY���易��ov�Ү�������7�vmu�ͩuv�'	*�$!�0QSN-Ai���`�!YЕ��oy�Q�۶��K@�k����s�B���Í�5�"brf%1�(V�v���d&�1���'6�,�[���yt
hs���#Pz�.�)���{�Ȅ���u*;*#Y�P�Ld����)T��28��Lgv�Y�a���܈F��h޶�Z1��/��k�Y����wH��[���,�>���o�:_�PnW�x�DGk�|\�]3���'�V�JCoEry�_h�`f�}�-��#F����(�K�c+�<09�s�.���VW)��P.]*m�h��{���"��!K�~6*�욮�:y��s��
*a�a>�%b+(ew�.�;(t*���9?�����OO���ez{6<ľ����6����:TR�/1b�O=I��̼O;�k�"��آ�����]����v�ﲌ�ҷ�n�6���86���������Me@�Z�ɦ���бNh� d��iq,*�ߟ�yac�aM�N�n��y>�(>e����E1�ҫy/�6��?/�9��-��.C:��lz ��
�$l�M�aڀ��؆�巈��,�e�|���A9�#0�2wϡ�~󹡚m��\�i�&���)� -w�������w�i�T��8貑��.�)�A$�Z��i�����p�s��s;Q5X�Zd�:?$��Q����fԵ(�I��i��g��Ƙ�0�So�oN��A�K%�^��"�;�Υ�[g�T/\rhfZ���@V�a��6	�t�|�zoYO�9ě��n�HKo�G�Lc�޼�p[@�6?Xf7�4�m��<�t���ʨ���BY���𠨝��yd5COP 0" N?�*D���Z��-ь�X��ɧ���=��������#d��Bf_�E����"1@���}��-Qã;�9�n�\X ȿ�{��c�E��a����МR���+���}Ә�}��M��TFn��D���g���"l��G� ����� i	6���y�C`+�b��bep�(7R�E�������@�o�`a7ݘX�1�k)xW��T��6��S@�Ȼ�xO2t��s����)�B�JD��꬚4�°�f{%�x\J�������oV纬�$�Ei�,z �w)͈F�v��w�Y��D�b������ʇr:���2��\h1���y!��	cn'��������8~bu{,uS*ډǂ�����-��x]����0"��퉯�ڹ[M�P����hf'z�t�L�?����֑w={�`��Å:Ӽ�����^���Ѥ������.��\ن'=�_h�RR�>Sf+Ƨ3Ϣ��ڰð�� aMA���U�e�TH�P�g���)q�tA�%]a����_��L� Y��AfyI����1��@ㄎv�M�I�&1�g�N�`�V��dyO�Yl�EZF�-�b��m��3EI��a�ō�Er��d�D)	�q}�/��;x�L����.���e���U�����2̤��a��y�)��ҨJ���,��d�XR�Sf�u�K	X�v���9��5L`;�$��KS��X�A��t�5�Cd����2� TG'���ŗp͹��u����CO 1�9���%_����P���hYJK(Kail�6/��!�����lZ���؂%f4\͌C�R���3���� ��kk���a���j���l�}C`�
��,Ӊ���)a� ��#��	�m�_�=�H�J�\��0s��w�
NֆS`�+t8vd�?� [���f]�
Vr���(����I��j����v�Z7\�� ��7�����"y��ҧ�V5����9H���:8Ou��`t�M��b��c�/I߂{�Lozf�&�^��n@K6lz�-Va�l-�p7�y'?WUJ!v��F����羸Y��:���I/ێ�۹u�ށE���I R"��U�؀Ҷ7b�{(Z_b�����3��y�#�BC�22׍����H�q�z���AE�eZ5wSk���P^QyD�r6�:�6�#��7��Tc���Z��ӤA1D���������L�V�^��E]wsڏd�%W���e[@5��	�3`����lb�"���zu�Ⱨ�I�!����"x����)~�8>����W_<��},u�N�ɴ����!+���a�����{�򍀂��	�-vIJю��γ`�$׈$�4C����U�*혿���lw,^�֣c
ԑ)l��9��i�	wz�����X��e��{�2Eb �����f|�xv| ��}
MuͰO��^�D���z H�ہ#h��t	M�:�`�c��@'>���q=�0*G���+��~�N�.=�RHSU7��Z� :u��eo�9/-��o�d6�=���m���MvZI��r�����SH&� _��䭧��s��9P�=���r�hl�槮w�������d�?Mv���;Tf�N����Ob��S�>&��Ln<��	��z��ѯ������M-:��E�]
f��c�0\���)e���^�jh�Y�9���U�#��;�-���zۈ. !����2�j1}�)���&tRNx����wxC���>�xw�O3�^��0?Z	��L��~�b��f@ �k���*�M1�T.���N�����΃Y�M�<gh�G�L+�HȃY0�����e�D��Op`3��?���'���G�61X�����&����_��U�IDO:����W�~ί�;	]#�%�xfMR���@F�r���a�ź[��q�����H� ����*굜嵯>�n�oEmr�'f��b}r�כ����*6l�x�^�Zr|J�EI�|�Z^����+A���N�s��O��������ך�r�C��ho|�њ/������Ӫ �9""�������فEI� ynw���R$(��c�V3+��7.	fq����A���k}��Bs����D(�~+z�`�Q��6�eG�j }��Gfv�~��{����dھ�����!�%�H��v�`EA��M�e�T*����+ș����2x��	���L:�,Z&=��M���=~rC;�G�},%Mt��Nr�"r�V:kn�.��@��� f{R��7 \���]j�DY{�L`}7�,�09�)�Q��7n�>�G���s�{�9�+�#΃ݦd{��Ij*���Q_���;YI��]�$H�5_#>I�bB����v�wǕ���)��m� ���6����k���v]�c�c� ��m��sݍ��A;��ą��Y��K�)pJ���#�G
ދ��j���9��Ë�n����M��x�'�\���$쁲�c��rqf�1w�ܭ?����O_�8��赱��?�_����ъ:��Y��`�-F�f�U/������ӌE�����Ě��e�M���WC�YTg?-IЕKT�s���Qы�a���e?������9aŚk)P��љ�����[D�ZO�΃�Y�@�r���V���G���b$#0 �$��A�<"�4�3��x����b����)4vA	�ҌXvfQc(���8Q�?y�_o��՚���4|��=��IoW��������HgT��묩�����=�)���x~��xXH�~�>0ɨ�Nu������x}8�׃�=. �(�^��\v�A?�2�l�3�㱃=����	�W�����DL#c}<�p� 7����v�;iY�L��kc�X��yh�x���	���}R��_"S���ˋy(S+Sjɗ��*:�\g�S�\��`��M�2�$c�|Z��ϫ{m��7Z��������V~dCz f,��&ׄQ����{�� �P�=�7,S����z����P����t��T���}IA�����P!����FdB�m!�"_E���,�>Y�0�Peye!ژMm���  �N�^ԉ5hv����ZcS�6i;#|A8���v�q���D~�ۓ��k?�D�0"'��NiU(bc
x*ɉr�"��@�iqHVX���E�_�k8:k��Ԡ՞Z�,L<�u�jW�Y_���߮N�S��n<���|��G��M^p��V�a��l��D�>>��ǎ��z'	ObHX�Z�G`���%�Y9$f�����g�|��uR�y��� ���5��2����g���RM=�}t4#
i/R�}Aq���k�ܣ����1�ǡ��4DM��a����}M�Z��v\��9�-�N�b%���EVZ����q�I���}s;0��wu��$4�疛K�­š\I/�]�$��J���3/xiX
5���2kB}��Y0�"� ��*�����(����-򏮫�:�����,�ޞ�p��r�jqW�P���o-|S����M�0�<`�?�ɚDRH�/yoV��O��+�GX�n�s��ȶ��*ʖ�>欒��Qk�O�
�.H�}r�\9���5����p
U�J>��N}LI���~�p�"[�U�d���țb(�C(@��#�]` �?uaF!tX1�Y7� ������s�@���4m&U@�TU��$X0�N�P'��`a��(��Dt�|f���c�{��n�q�q�u�ɾ0��f=�`i�_��*��S����%^����2�u��	�{"4}�;d	������f��c�@*k󘹐iO*��[-�J��P����,���U/Y$��ND8^�쫦���<��pC��S�|�VbL�Wΰ�eZ�g#�BGC�)U�i8L�~^Q�6=!����1?�u�p�t��d�dZ��_���|,������h�Ǎ��9����:�O�1�O-7����
-��Qf�uU;�"�g��7�e�zC�݈C��Aj��MiJ�S�zaX�p��z�1)΅2 >���Y��ѝfE�Ic"��I�s���2�׈�!�:t(��k����ڜ]_��	�h�+�S>�E���T�$�Qm�%z�	C��%ؙ<�&J�z�G�04G�0�ҏ�R[��XR����JQo�ǔ�o��%�9n�)�M�TK��2�/ ��7a/�aջ�UG0���8>L��|�e/�]gf�!��i �aӤ����`�������b<���=������FƮ�js�Ւ�d�)�.���d5�*�Q{�}`
rϕ���'�댜��X�X�p�q��P 1Ew��B�ѪWV=,���D<�P�f�p�P_� 9���,;/v��)�މe���<�ݒ���;���1nc�VD�f���aA�d?<�}�EX�����7̨�e6���X�f�?��n�O���Qc�>e':�����]5��r�8z���XG�Y�Ǝ��G��]��y!���8Usy��+(�u�oq?n
�
�f�Bupޗ�78f�y���Iq��G:כ������������z����[����3V(���V���g ����	j�Vl����'�"p���ݵ�,"�������� �-�뇥��g�88iٕ)�M'�:$UsX--`���N}<@@cjk
�U�y1]}5SrI�;�)������M_/h�]G\,:p�C|�h�a�����[��/�O�-7�b�����o�[�/M�	��~�o�w��,�@�w=��i�JM�m$���J����;��="jU"�<2v����`ǀ�z�C����A^Y@Kxr��Q��21q�"w:x�������#.���A8u��1��ū|����>�C�Ϥ���`����(7?2 ��C;��ZG$l�����pD*�,��-d^^�=��/�G0DČG;�hl�\��󻗜y������j����,�y�>yI��6�8|������]�1����iwp9ˁ
�!(d�ҧ�tv��	�{׍��w@$�]y4Tdo��D�����z/8!0�,�����9�P1?��҇�ۧk�Wm�1�Ox��wІ~?��G\�$��]^]�o.µ7(��֋�´\>�o�6���oݏ�'��f6��\��jFw}��ФHx�����;�p����p��E�T��X� f/cg�
פV�x�`V����	|���A
?��.���5\9Sh�ю����:tk�Y0��8<Aѧ�6��Di�9�S�������eF��&Ćcƛ��7�R�K�nqG�]�
R�S� ��?3�, �ק������LQMmZrz.4��|뚶�C�D����%Fp��dݿ����z�e<��4����:@ā�2{6�㴫��@ Z�r~pd�b�=s��.�!�:�Qп�˅)0�ۜ�3��v^;�5�kN
ɕ�[I#�<�� r�k1H��n��H��3r�f�O�)p�|��
{��p�����]"�����:�2��Z�d��niHw.W���Z��Y�5�'��|��؄�M���W4C�CK����C��F54ˆ'ĉ��9F|�P6 AZ|M�'��3�J�{G��(��xE�!%�ot;�Lsȉd�9�j��g��%�H�ޠ�G-W�GBdy������|Mo�p&�<֎��>5�f�>�)�o�Xz�� ������Aw�W����hvWs��Q�FT����U�	7�+�`�]s?~D�N^I��͊�*�Ɖ��)�qRya�|_�+0��a������X�>&�P �t��^��6O�M��ޢ߰����=�����ᘮ�S�2-�
�7G_>�v�,z`#��!U~KӪ_��Rw	�� P��ȮyO(�_	����f��А4��$�}3�T���#�X�����D��żvT�хi�J-�A	�kY�ꋼ��Q�V.�P5$�j ������hu��Z�K�܊��SC��f�ꃱ�ܬ	���#��2��+Us��38|=��A�$��{o�YrNG>b����%�yw�m�;f�����5�Oj=�[v#�a��3���p� 	y�-d�l=&�\pF�I����n�vr\`�XK���={�}3���f�p�q�e���[��΢�J�M���a_^<�<�r��y Z�-&�{���pɫ�{RZ��?UG��2\�,-d�4�p�&�������Vk�>��9jW�-kxY"�(� ܘkm�أ�?p��su �lu�2,L���;*;p=�;���~���9�C�sB�S�����i���&��PB��q� �{�c�T ��O����S���;������MTJ�vE"��h<Y[8g;�h�t�E�߹g���"G�s@�:���'��H����7g^��^���m��Ŋe�h���Z(s���g����j���� ����Gj�?�X�*x�d�q[~a,��6���:�/sԲ�9 ���V�(����:$�v\����i��$��Ya�B�ڽ�"��nzhnmA������TZ�g���p<��dT��~�T�ޏ�����%�E[p�_�Tc
w���WEY�wqd����<\'
��|�!y��������,��w���E(���gN�+'T%�1D����FC������c����6B�Yz^��M��� ��h�u3�����B����}bD�����7��(Wm+��!��M%Ӝ���^�^oB�ԠC��g'�o� V��������S���� ��ғ���<K�C�(%ގ�d��$k�B�l��A��,�`��r�ic�zx��jg���J`�Ѣ��"�?7"Q$o�=�@���_bjO`L�x��b髍	��s��a��zA�
� 
Mb��u/���L/�$��]��Rws>�-ܰ^���u8��L,��R�ۂC�ʏ1wyNDt,�`��t1���	���E�]9�i~8T���b��\���0�C2��Č��s|b�i���w���F2����f��f�����*��/�!d�Л>�Z����0��6ԃ�3� 1M6�]ZY�^}����jw6h�d�jԼg��ZS�@m�Q�Fbw2l�*O����^`���bmz�s���3[ �UH� d�z��I���{A+�aX�eh����=3��x$��!���,�R���b�u�8�+(L�עǗ����'�=�d®@w^��to�RC��Z����R��z�N�5��y�\J)c<	�����f�<c�*n\=�0>7]����hXu����ɮŹLm2 ��;���稤���z�/�S�z�W��o5��y�-utg��%�hJZ�n1��U�gT^��8�B��I����Vu3�״���"�{�����!��|���,䥨�b�Y=jz�[Q��*�&eu�Sdo4��*s�7A[��o�ۇ�I��ˍ`��yԼ~<2.|�C��e�0c����9r!��vj�Mz�VX����
���w1W u}߰#X��)�1������U����HEQ�0H>չ~jc�C�Fϵ(&B�U�E4y�Gxr�6<X��j���H�P�K�V�	An�LkJ��>n!"yO4�݈�_䯫�A�t�!�z6���@Q����Q�>��&,�t�!����8p�l���)��7�\����Ag�l�[�6ΰ�?a3с��jᚇ��-���ES�[	Ś>��˯�Ɋ5�9��4��N��R���1�96�WI宇��3Rdh�ҨʜJ>Jh{-��j�y��K��[�Pb� D.'��3�(s����z;�2u��j�me���S����p�ˎOz�(�S�� J�Is8=�u�pB��)���se�7�y�<x�ef�j�*lE�2�
g_5��?%������v��f"'I>�Ɵ�1����lU���<���2^� ��a-����R�R�eK�'����L%�T��`��� ���gL2A�M�׍���1�y
�ۿ�B3�ʟ�xq��n���Ȅ�*s����6����۟���K 0�����5!���͟�v��D���Z�����;�$�^�<NɀXs����Ϧ������j�}�̝������*{��Ƅ()���]@n�
9��N���v3�M�0VK��DY
.���pUS�	�wV�f�7N��V�BMz�ŢI���c��Gӿ���I^���]�|-�uf\w��	�Y���RF��Y�+����qS�nS�F3���C@�@?�g����u�h=�b�*_흀_��޽�e��we����1s������2۪�-�3��Y���@�c<h+�5�L�A�d�8�t!�I�k�q�����«O�f���J��ɉt�E��X$��c�Z�)9���ҹ��,�=^�V�b��Q�#�Lɟ�er[��*G�T�#@��`j�M֭	����Ԛ�bՂG��+v"�E0EQ��
O�BZ$K]W[
�]k��	�8`�����TZ*&�H�6"�\����?���Q���W�¢��w^J;q��97Ϋ��۽q��k�L����>k'�Y�Z�@A��i��ȩk\�{r'8��hm������i�����c�$O��?��{��+��]�C	X�IK��r�; 6�M����[�e.P�E������\Y*b!u��İ�,��J�;G�n�f�8D%dO��t
�T��'���]�8o)X&�i�жM���O�޺���I��0Zυe8Mr;��J�sFDg��P�!ɇⵆ��!ëHr_zX�N�K��=)Ʃo �^����ˢ��Fѝ'Qgw�1oG3��3QW�{T�-	��"��q��P?�ͷW��6��wx	��S���?}wU�D6o<���7�/�[WȜ
�:�{�~��*�Փ�g�&棷6r�|��-����dx}c�m�F��k�,�,�{��H�4ӕF-~l j�4t�� ���Đ�J��f���9�gC�MթX��(~F��-	��4����U�G����~�f��P�C���"�xN�?3�ʌeVm����l.~�BJ!�|,����b13:
]1[�;=�A�3-���AnD��mͤ�ܢ��?��A>�"v�@Y�1o-����
G��ܸ�+��x^/ș�s�J��Vz���h4u����"d�� XW���q_p��Ǥ�7(9�6J�Y�[U<��Iw1dT�[G����M��;%��� �fM(�����R��������A�8}+������X{'��L��ć�k@��ŁG�`�\4E��Z(��������4������rih���Y�])�ԝ�-���Qp����>��i�sw�]46oi_v��ƘF��L=^"�G�+���y��������.	�@��q ��v���R�pe�7e�e��tէ{p<��4��
�_����E2}�����L#h�{&��|9�U	0��J ��3�#uPA�_Iu�����������Q����������o��g�>g~C��sz�r2�@��hIW'\���t�����~�G*
��DPh?�f܃m�MI�umᎲd ~�90�|1��Ҧ�	-6o]a����1�
�a�gx��s�c-�,`�l�is�g�-�&��ě�����=�3���hr��z�f�ؐ����^���� �څ�����=I;��.Y�e����c����`�O������Mr7�wy�N���ڋ2�^@S�ɷ��l+l%LQbS�u��`%1�6
��+h�g�S#�h�)�JJ&�@P�5���P��3���h�H����k{��_��Cz��vH
��/��>M� �B}3����[@1kk5��>@&���;�W:�9�T�$���~M
>t���rq���:߳;�1]O��Ͼ©�����D�	����=B����"��º�6?r��diU�  ޤ?�uI�{���4ŮQ������	&�1������ ӛ�����	�|��"�n7�ͧ��g�Ϙ�����vj#F�O�@���gWZǈ�������U#���&,��-�2F`\5ؐi71��s;n=�,5i���z��������q�l��W�������ϰ��i�!�i0mɲ�J�jIˤ���m����O:��OA�nHý[@���;�z�E�Qq�^Ȧ"��+u�����*n8�1�P�إ���(rRfa��-�KX�M~y�|���m�	����#"VÒ>��i�S]U*�ᛝ����4I?����������%r/�����k��8U�S�g��x�ek*�"��#��p�d��1jfF������KhG�C�*}s:!Pߟ�ٱ��K)�f+��&Z�m��⚱�ѯ�p(�R�n?�t���~8Q��<��
�D ��-J�
�b�0��f��g���"!ФՑ��B����B����͟2]]��{����O��}p^J�p���u�D@�a��*i<8|�9�����08���7���ΘDf��c̺����WJݕ�x�S��k'h��ǆ�"�uO�:2dw��
\��
&\"����E)���gt|�}�}�U�z� �s�)u�/�c�Q�!8�C�Cwz������u�}G���1bmS�=����1"EaFf��Y�����3Z�iu��Ѡ��]p�8��ñ�ex�H,_C
R��������ԷZ|�4ޯ�[��EO)�6x����3�3j;�T�����RdEx�q��k�.\
��u��#ι���2�s�l��l+vL��{F��>V�I���%�TT��ѽ�6#o��Pe-��>UY�=G#�ݮn'����l�2`0��.;�_z�rU�*;=6欈�^i��;�6�cZ9�y���+ф���-�>�a@[HXSC�V�BnQ��b���~
l��))� 5d���N��=G���WU�eкP����O �Վ��^�b�*��m��ʏ������	1�3��{5cE� �n��M�<��(o����9B�Gli�`ɺ?3W�m���V-����J6!�����h����8\�6W@�UL�g�}�{%��� q�┚PrH��/�]ߎ�3g{\d���.�����Am%��~����&w%�<���&��)���N�]�ŗ�"�M����9��⇡��\q;T���Q�Í�mk�L�R�J��4}G�%��L�.�y}M����c�D�cյ�W�r��s�������xK?�}*=��k��($UG�Bb�������&��F>_o��ۅ�u���C܎���>$V6��a��M���=^�Z�<��o���8�>ݳ>�/���/U�}x�LQ���F+���i���e^��Gq����.�����͟ǎo�5g��K,?���V+�O�cN{Ѵ��=��xq�t�ǘ�;hÒ��6���j�m�
�Հ���2r{�}FO�,!ՆG��Z�Ef5�� ?NВ6�:n��ol~��F=�����Ek���1� z�I�}��X�~zS~�Ï	�Ej�
?%#�$��u;�a2���k�H|�v��@Ԋn$K��@-�|���WL��_�K�Sx��2oc��0Kz�_��Oc�b5��Y��b@	��c^]��H(]��K�p�&�Ey�g׍��Bٙ_`��Ѳ&'8��H�tm��Z>Z;���$��b'%k�t8�g��b�u"p7���ޗpjk}ו�ĥXXc�}pg�<���G��S�5��d���e�Fi���̲5o䔐썾]���5�%7���J���M����.�U��G:v�ww��B�6������ĞR���؊}��u��¸|E�j+�gc�Zz�<>tI/�R�6ϛ.<�)�Τ�$�
щ��.�§3M��������^4���Cy�v2/Bfc��ф?zf�U&��_7�)� wM�p�=4�o�|8Νn尰�I��ZM�����!F�?62���sD�O50BR��X���� Id�#��E�c�Io��^����!H�+���h	��~(^��J�����,!�Տt[�d���N�5!m�r��;7����I��@�,.�l)�����q��$�f�a��(B�t�_��T/��8��V�[	t��r��fn�s2�W�V�LV�!=��Hu�I��-�������\O�!����6h�u�&����2�/�Z�x.���A�ߓ��Сh
Z�iZ�l��t� �a��K�I����Q�<
8���p"��R է��a�Y���z�����d��4��(�K��^H� ��x���1����U���j\�����ʶ��^7M
��W^C�7�)?�iƉJ�|g[�[��oŊ�Ȗp���Z0qr`��B��$�����9��V�;�p��P�L֛}�W���|�`���w4��7�Aߤ��[�m��ǵ6���N<�"����ׅ�n~�ܸpAG�����쌻��ż���YTص���>O5?�rD��P��+Xg�-�g����dU��U���C�S�.�3����#(�E�'�F��l��J�Y����`�eс�v2ŭ^�� ���A��:��tܟGЀ�=^?	�蕧V���]/���yD�;��Z��=�$Q�)��Ï�͊���	*��\K�8q�qDȰ$���F���s̭&����2zf�&$�����JJ_œ@B[�񂇊�Z����hj/�O��i�[�2;�T��0�l��E�+N;s�#
vr4hI����IJ�l\�6R�����6$�9�ۀ���g�k���Mcm��f�
����B_�� �������r�D�-5����E��f�$�1!�t�6����Foy5&�ew�Ԁ�]�Bɀ����Krl>১2���6�!�_����f�������>:9Љ��{^���	�!;����^[���1�G���`O/�������\��Z���K��WP��|��/�,h�ڂ~;85���-���pN��Sz��
�yWs4߽�6O9��|1�C�NI�۴�,� �t��Z��A���%���CyUH\fݷ.W�m�(D˽}�
>Jf/0ET5h����O�=qf.*FB�H�ŧYv6�U]��I��o��r����]��(j~6G3�.]\O�ŧb���0�D�f�x䲟+{^��n���f(�l0gzC�P��=�Ѻ��ͯ�pߋ)`(��
xU
i��Xzi��%X�'����z�D��h�5��TZ��/�F|��U���jN+nt9��=a:5_ʸ���\�b٢�Dv�umN�G�������f��/�m��I���]�	�"�k��oJmh[g�gK>�T�.�'w(�~m]S���t�C)} P�]�8�482.�*�|ݧr*�������Hɟ��ҡb��H( '��o���t��&��]��<G�������F؟�����c����WZ��N~JK����/�<���?S������E@��N��c�ܧ����� ��*�wt����T��=V�UJnj}�>|�5y�N���$�N j�p���IT��ߤ=-YFV`�P[�Z݆�o/pv�?�u�����ȕx��]��SP͓K���1l����5��倩k�n �^D�hF3��i���̬�GZ����3x���8^�����
*���kZE�?,�[�m&����#W������7)x�}�ܦ�]+m&��q�M����ۺ\;=�ܡ�_�-es,������ea���BЋ��(@1������S�@�3.�/�ȗ�+�{kYzr��ďY�Nz�wQN`��@�!$F����O���j!`�P�@"PL ������l��MO��r������4�x�(�
�2��%Y�wj0��8.ќA��;��_�ca�c;�.�3��m�j�ȯ�ƪ�R�0<�� 3��-WB�rȓ�N��B�|*�o%{�y��=7���}y�k:�lK4G�ۃQ�6�㿷<�J�y��4����Gu�͘Y���R<�8kvR�\�����b���l#&2!+��9��[��L՗1�O��KJ�P���xp��O�ޠ�Ӷ�kv���_^_���k̮j��݈?�H/;��S�F��0�e�dm�A~�ئ��
��X�?�#.�@��N�3�}m-�f���\����6�Nލ�4��9lP�ʰʖ-dɁe�ń����ss�i��
I�
l2�?�C�T����4�s��?F�q��Hj�m����K�H�簭�n���G��P����>϶�  "�m�������֜Fꖀ<e\��s��
H�/m�7� Si�b�޲7q^�r�D����x(e8mb<sxn�U]o|R_��.�!��#Pds{�"�Ad-�rh�4~l@�T��Qe��,([ڢ�~\��|xu5j�,D	��x ��<���f-v|S&��MX����"W��r��@�Yܺ�/c���N(y˹_z>��١6��Kd=9i�"tx@� B�O���'�ث��m"]��T��u�vB�a�CW�띥�
��wE��=o���n�E��Z������y=�K��8�c��I�(_�!HfA���4�v}��̥�!�,�8��*b�9-�v�<	�/���h���.�=�0�fNE�}��{O@��E��sXm�\(r�g4��j�����AX)AB�ݱ�VI�t�����)�8�y��4���`�������]�M:�
�'U]���_C��E��.��4�C҉@�)�%�� O<�P�:�/M?������>�kx��x���Oۂ�Lvǖy�3��q7��#����T�K���#���#ŉ�!B�(�ŽY
l4!��w��51�Rä��_�����[�6Y2Ŵ&�N� �u;}�P ���0N~�����.�Eh.�Yw� �_��#�׻���3�q9�fdyU����7&�C�6*���i0�Z���k|JÏ�B�xap7��L��Ԙ(�ڷz��(s3B���5m�T{�pj'�vv����F�ɬ�������l�_�ҡ)=9��wt��m�|�|�+��`��ʐ�z�b��44K@�1�t�!�q2�z�6���A����U⥿oʂ~����q�J�\d^o�^pJ�
�}����f��\Ymb��8��fC�Rv���y,tĊ�Z!i6o�e"ho�����h�O1�w9t�hL�����)&�ŭv�ѷ��2�t�vE:[#Y�A�0r;�����
�.~���S�X�{�z�$n���OX�c%n��1$��]OO���vzF�Qՠ-�2<��`���IJ$�����A�2m�yn�֚`�I�����Y�tm.�_r/R�8�HB	���~wQ�F�dA�7/������!Xf��X�U����&�;]�-�K�lQ�>�Ek�O�	������l&b�Q:xP,�_jg ��,6�f�.(.��m!�&h��@��E��W��z` ��k��Q��תJ�S9pm��K4�n5��~[g��W/���B�1��_��d�v�C�Bm,9[V�P< FJ@��h4��훧V�