��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�nU%��l�F�y��7�R9e7���}��3�)Nп?�j?+ t2���|��T�Y����œ~�F/���E��s�		�}ѳ�a����r3m�X���j��DT��bO{��6�t�#v���`�&�54��Q��bN��I�![U�B�,]�w�r��b���b	 ���5��G��r>��T�CF�I�&������y�C�)��QNF����4��'Qj�x_`�'օͰ�x\�����~�;��˄lB����8�Ѳ�RNrB&���uS���o��w�!|
:ϻ��G'S��.��Hk��+*��Y�wE�*+ ��^�9W�+J�k�ױG��u�� ö�L|yO�K���p�4;+���6�ҥ�T\*�h��9�����wg��p��Ղ��,���Գ�m������J������]����m�[�ۋ˨�5!�ý9?X�W�x�Y0&�g�Q7�W�n���3�a�3{�_u�or\~
��h��#����\Gf�7����O�8-;��E��V@~A|0q/��oѨ��p.W�HQ�����" 9 ��n���6�;��&�zb`IQ�X�Fuv�c4�>zK.K�|ZFz��ڮ��Ȧw7���t�=����?q ������m����s�*�XR�����V"�Q�Б6"��|���Rg�sb���P�!��D$}i����p��gQ�!Bj#��7�h�ch�����*�{�%��v��b�rk�����#CE�󂉢W9���)��|�K����?p0��&�~4���T���t�څjc�7�v �������ꯢW��UjLx���=��S��A�u�pkqs����v �F��&�RW����<J$�&<X/��R+��nn�t!b�D7"�M�ׂpA�5���N�U�ҋ=ͳT�]c!:�c�dI)��3F`&������x��9�U"��=5Ka�P,�X�b���4='xq�54�~�.��3�,~I�tRl�����R]g�@�N����R��v�qD+|<u�2�"��h��_��2��(Ry2��ܿΰ,��:�D�b��T�����G\5�ض��|0��N-3[�%:�'jaU�n~Cd����mF�t���EA+&I�����a�M��C�ǐ�Dg�8�b^�\:�NfR�w���c��0��e*�14o���*��f���(o&Qm�g�~����o~`���g_6U#�e%$X f�Dlի���
��Ћ��8���s�Fţ�6����՘W��&
�,�m⢐�k�
ZA��\LuW���Y@Ə�93�E`J�O���3Mf��z���ۋ�ўh�m�v�b�v�7�8y����@�G�2VG��U;�����R�V��s�+���[�Ab�(
_l�څ�gˑ�(��GQҊaU�6�tOR_���e/q�a�5[~-'i��<^.=����q�\�}�T�p�\t)g>�C6�֌Yy�N�0|�wK� ;����ړ�=H>����)z���6� ��6�V�_z�Y��r��8L��UWM�	
�%84�)e�;��E���G��G�zd�&x��n.�Y
ˌ�s�rЋ�����Tyc+D�GR2���Jz|�� Ey�Zј�a�`5_Q�$�#�B�y��ʼ$6���[s�5b�71��<"�����/Pi8ɥ�;Se�D*�܅��L��=OҔM��; i��ʒ���KFHl������"Ǐ,ˊR��f��s��SOaf�7
{�@���!Pf=����n�м��&�y� ^E@��.�a�"�W�%{i�i��jaJ?��c�*_�{�ܱ�I߰B���l���F��c-ĸ2m2	���+|a+k�w�)���A�w�A����-��]���lw*1�|"Na�!�����@G��|��)V���;��r����;�;E�����HѤ	$?;顾���y��jA��9{��H����·�Q�(��o��u7�VY|�n�νpWW���f��R�Y^GǛǋ��9E�]��8t\W�j����3��&lƛ�os��m[�L����81y�ut{*�h%����_�q��p��4m�0�f-jiT#\=̅��u
Oj3�C����jQ�*+�)�ul/���x_T����a�z�y�҃�����)�	8���18���p�r$�ր�e�dbXDը#���Mx�}�bLw�rt�W4^�"�(�u z�����8�,d��A�-�LCt�A�W�y�ۜY�|�xd�ִ�7�~�BN��ko4�0܏|x8��V�H@XP��+&�C}a����X��v]����	b�;� �l״�P̓�؉p�Y��ݖ�<��eqn����Qe�fH����9�\�&j4�Zp|i��V� 
�jx >TԆ?��B��nIg`��rwO��MTy@1@��B��k˅i�5j � �0��a�Dy�m&dGt��0�-;?*�Etu��]��~��u�(tX5�)�r��^�I��s-f����M�dS��Tx����F4�n�)�N��0n�[.���G���4�]'uۯt�����m[����*O,
|����F��| w��tV������13V<eH{q�TDl&�g�uRU�WH������}����c��C�]��������p��nn������k�ª8�
i!U �<p��%�a�c}�'�i(K�s��c'j��\�i�n���2��Wh�	=2��}�J�.�1Ety�ׁs���I`�F��yǾ��	첟���'L�a	�Co|��C�Ost�Q8��L�����ZC���Q���B��L)S7���G��{�2jQm;P_fW��ujf�%���Yd���iJy�Q��QP��E��*��i�gRj��	�b��n�a�N���]��;�3.]@�m��`?�Ě{�u��-o>	5;ە$��h!uڟ��F[��L���g��kIݒT�Mg����[��R������*����zbX�^�Ş��m6��ɭ�V��<x�V�/V)�T��Ԑ�1�-m���)��_����}����I-�ܺ՚�"Z��c��n���i�TxH�3z�p\E��@�z��W�e�����H8�c���O�������D�wV�Ĉ�1l�z �Y�
ʴ�ip$��E���H���,b�Xy��h��_����M���t�/��|��r�!����]S�k�P���L ��@�lʹ��m�����+IY����k�%��dkZ�L=��3���!Þ<I=�5l�G��k�Ny:],6��}jҿ��1�����H���1��#p.2�����!lڄ	��Ϧ����}����xv�֮���{�lN9*WXl�p��JepDF���ug�I���@��zZ��M`�؍n��K��(9'�� ��%���c�P�gSN��:�g#D�∼�h��44������ed葱�)�]��S�LX��7eg���b����O����/�3�B��>[r�Q6�r���R�����{�O��p��&W�&�]��w��i�hIS��euKo�{�N6|�eFʠ�7��?�|���^���M�ɀ��@�g�I|���r>O�|1�,W� �!�c
�-�f;<о��/HBa���]�(�S�Cy����c��u3J�G��~�h���/��5RGS��]W� �Y�����2��DE\�����S5����|��e��ֆ���4x�]brl[UW�PK��9e\vy5�[�'�@1�
�G��_9�"��;�p�4��F��Ee�K�Qlw���Lأ�{���V��g#߈ �`��͢g�f�c/����haj���cv����R!��y�azn��PSh�����SWPK$���Xz��c�66$����hT�SSF�P��=RxI�R(��1M���k�!�"�۸���,|�cm׷U}�[��#	K��!J�R[2h8Ƹ@�/S����������WHz\�S�)	N'��
���>A�a8�<�:����-��DE`�pú���b��2{~$������ �f©.�˒:���1VDoX�����0�Mn\fߔwK}�t�|y��|\ l�: ;��U������Y�;��@R
�ǲ!���o�?�n��P����C�-zM ��@� �o5�Ѵ���X�B4�q�$1s��q ^w�����N�C�mG��R\�mN���A��6~���w���Kע�W	�����[O�����(R���*Sy��@�J��k�u8X�R�k?�G�A����Kۖ�[�L[I��ޛu�D�#C�'uK�.=�j�eLL,^�`�z������_���2[�K���a�3�N3�;*��h*���D�_n��i���$�h�=����J�:��ZA��#��2(��.uS|�|>�4�
X���ż,N�#[Q��I��*,H7
�mHe$�:���p���;`��u3M�C��^��~#�	��ƥ{-?g`2I���5���q��!!���@�2^�/"��0pZB�1���T����:���f��1V`ʜ�?�p��c׏�
֮����UR�$��+|���P�:�,���4v D��"�+ŉqq�?�uqYpC��:>��( k�F����{�GͶ�=n�������ch�x�n�~-��
.#u���@h�L�h�!��?�am�;�I'4�f��vmRr|2t$,�It���Nv�V@����c� >�C�u��EwnC8=WeV�B��6VS<οꧭ�Ē�7~#��_N����FAݩå4]�5�p�CR�k���1�~�u"T��_�J�S�Y���o�$h���A�S;��<;eT!��5���7�҉͍�v$V>�����<��\�sY���io�B@�uio�kR|��-��p0�r�E��Ԃ��yx�G`sf�.+Ha��
2��h����Q�k�~O�ǅd%����I�_�o�2�U�������	�+���yv�\�t��+�,sZ0;��pU{c�	.�P���y~+�e��5#υ�Q髽�UI��6[��Œ�wEaD�;t<��>����V���k#�r���c-XP��M\��tR�3�KpR��� �}��P��]��=�Zl��t�o�	�Q3�����'�]+MM��4A�t8��)J�������)W��F�����}n9�1?�@&AQ*]'�������&���{W�#�;��:���A��h~ �>�"i2ѭI��/�:�6ocS���eW�d�Գ{0�pi�rQ��s#�Ų���)f�2��R�	e�%G	󀣬!�.d���4�|�Di�҆��8��e�Ů��Ƈ&p�W�^�z� ����2�����3I1���h]B�}5�8C5&��-�/��0��V�dJ�!'��T�1��FI��K]��?7V3����P�-����>�e86P�r��<�,In�χ|vS�5��ʀ^J
�j�>U����q�A4��)s.>T�N�S��
N�1TƭT�A�O���R��6dO�풿5D��YW!1��#b�4ڌ6_E�v��Y�����G��,ٺ�p������� &^t,B2��<����,���E	����.�c��Ѳ���9e��h��h����գ��'����͏A�C�.{�8�Ҙ�	\.ɃG/ŧ������X�V�fG�[��:�t�/1wp�	��y�F�0y˦����\Vʌ�U?i���I�M9QL�ʵ�P�=�e�����܌��׍����S�ܣrI���pe�:`!����G���@f�Q;av2s`;�`�\�+7X����+,�G�4��݁[*`���\7��ZɍO����}��m�ޛGlx�D)K$�� ��|B{�~�1�X��@`"x��p>ɡB��Ыl�n~ ���P�eDC�g���)��
�v��Q⫊��5](u�3_�E@���	���!UfFug�c(Wv]���rv�SU�g �b���s�P1l�3�x$Z�+.�ުJݲ��N������9)�4��<B��/����St8rOCNd��>�T!W��B��l f��Fi1Y���,z/�}frPm�S��@������B�@+�Ѱ&_��^�Ɗ�\��u0=o�.;ZA ��,��8�4����ff}�Oj$]��q0���R=غ��~7N���{ؑ�F��(�3�ޖ���W�����]r����Qm�$���bNI��hۅf�/g�S��� �,�.����L��|[q�~�W���]��9g܃�%+��c��f��rv���B�Ѱ�P�F������E8�a��S{�Z錙��q_~D�/䍇L�A�R΍cvp�lM�s���ـ���B�2zRJ{���2���9C@�e����m�tԲ�1���e���^V�	R.�W��Ϧlb>K8"4���h�}�/�T=�l����(��Y)L����]�P]ֱ���R�Ӷhy�S�(4,�?��bo���j�S~t���}�")fpϴ��|�]�]��������,ˍ��f�kr�5(��$�~gv6��.����N�i2�&R݀�����df+����k�;�c�0l݃�8ʾ<�T�ԡ�+C�!���ڽ<�G
u�Ы�Ak��,���ax�\�������ķq�
�M"���*�r�y�$Ъ�˞��k�<\�.8��s1x)�Ur�������n4RH�bx��@�v��ֺi_D�{&z����+����፭�s�5�Ͱ�n�d�w�V\���U�Oi�e�t\��t���f���n�?�as~Ըz�Տ�P��񹽌�=iehI�7[[�!7#Q ����S������Rg�I��aV�W�>�9V(KvӚ�����c�1�+D���D��t4D�����1K�<�美4����Q�gm�f�	�7�Y�[��d#��0xK$��+���Q�u�Ě�<�҉}����U5NW��o�LWDK���c�vN�U�W�R���9�����������c+���/ɵ�W�Q�#ht���b�e�
�0��hr�Â�[w�2:���r*U.Lf\b��!������gOi	A��9����rcZ-D�o�l�:i%�YC��0����}�7q��؏ES��G�ΠI�����~{�e�Ӧ���:�B!y\�s0������^\ ?�&�u��`��r���	eJM�KK ��1Pi�i�������Y�gI�1D�
!�g˞����X��.;��x_�Pp�aay����w���[�K{#����E`��� �Dׁc}���t>
�E����Vz%C׸����u�����W5��{{C~wi[�{\�K��%j�m1�g��X[<9�أ��|�#�a��{��`�~�.���`V}��5qS���Bt],�[ �H	�#���{�>��>�ل���׬�w�M5-���b���^���_ǫֵ�F��f�S�(�.|��h�c���ڞ�9��ڹ(�.B���מ8���6�Wz��,���X7g��xW2
y�(���D���M�����36�!�g"A>ޘ�3Ϥ����pXT�Q���EF� P�f@UH�5(�f�2��'Ƶ���w��Y�ɑ�(�=!���`�`�Vv)7r��I��*Վ˃�Z�muN��Q�(g>zƿb�4=Dg�:� J[jq]���wv>��_�z��o���Љ/"AL���Z��$ƕ!b�7Z��;+N�q|O�E[��p~ɥ�>���aTe����҈t0�a�Jw/�m�Q@��A�ľ_.���y���j�6���2*��#G��Y��g��2��Ԉ����5[H+��$%��E]kF�s<K�����-��%XdV�i5v�Wü��ب�Y9&l���A�q<^�"���ɇZ�o7����0Q���Hy#�^����r>�|�s�����԰Ҁ�,`Uw����8XR��`�QИs��%�Fa-/���E� ����x�B�fp0��X�NCR�Vq�Bbi���v,�]d��T4KO�z9uI`�R�1��7S�IS�/���W����fa�3�d�P��9g�����I:�X�S%^Έ+�/4�캛$s�o���Z�[$@���~�2D�n#s�)�P�;����>kw����xp�m6��y62;3�H&,�V��%���{�0��%�����8m�	�^�hP�b�J�_���K{X)C�(�Dy
a�6�kC 6l˔���nă���x�PP�c䆂�o<X!e+%�X3[����S�dP���Z�Cr'��^�N��!!��Dh�C1�#�w�܌D}jO��)8����C` Ҍ�^-�x��i�[���Ϣ�1��I`��B۔�0Z��2��/ܴlvɪ�]�`�����w>�;[E��l�(�|��Z�z��� �㌞W����E����X!�$�}������d��g	��{�κ��ʟJ��r���*G�z᎐z�T�xhkkq����X�q�U�zL.����Fl����nQ�q*f��yj�$2�y�7�R;ݒ��:]�X1(��s�:����#�����ۧ��Bp��Zr7GoB�$�������k���.�!�S��O�טͼ?�'S��R���q!?֞O[ȝ�ͷv��l]Sޟ 1Ƙ�8��MA��Wѭo�F�"D|��Q>a���\�mb&K��X���F2S����$��������EO��x��&W�����[� �(�VY��NP�c�պ�S�w(~���8�N��������,T��5`u�D�a%����T���J^��3�}H֣�����`�<�Sz��S�+9��DR�e��G���F��/
+�9hA�����g�Z$�L��i	.s�l㕅IT �d�|!0�Q���q��0bJ���Qx���4Ψ�zy��n-A��W~�M��TV�|���)z��JO��5i���C\x0OL�#G��h�(}J�O=JN�xpY����)���A$� �v�s�UcdDGB��6�����Dx�{��w'ifj�U6h:�s������Ty_ d�	(�y��V(}�E�1d#�R�}Է�й�?R��X�2�)�5�iaD
��]��l�Uel��1a����Zy��\��J��G��֒�U78[!Ȕ�;#D��M��3��|r��DxŤفܸ��NB~�]O{�8lͿ}h��Dɏ�B��ܴóa�~�����ysuQ���a�~k���g�Ǵ��)�+�Ł��q)���I$/��W�쫥ؒ<l��L�K"���c$������� � B-s!N��k��2L���>��C�}W!ۀH�mNh�b �=�������ݐ+j�����=��j�[����|�Z~�CB��-!�)��{�%C1x����jo�� ���=.��R�9h��!���©���~N����8�g�U���Յy�H�HR���B�3X����C��r���"��,Đ[���6���\��G�v�*�Yu�� Pa�I� EV�o˹�/-}Lz���(Ҽmd��XEQ�l%��8��B�	��0��c�HpX������q�ݍ��螽�$Pe�Xb4�X��i���4>u�/���+�C�X<Y�~h�.T($?�Ʋ��~|�a��E ���)�m^I8��zp>���+EA��y��^}��2Ag_���|r\q�ux��;��B.��z��8I�CX��G)�H��S+����ǂ ����cm�.6M��bx�|.���%Fʍ��_Y�[��t)�@�d�o5k��7=1gU�^�m_�ٸ�<>8㖡w�9��k�G}�+�V��[>���L�6�
FN/)������:���qQd��]����Շ;�K�G$�*�7}�\R[�kk -����5v�(�F����X����E�5D�l��#/m�}���� KsAK	���v}��)������6hU��~"�<z��̸��V���5��=B��۔k��z���h��к��C$A����,N8�d'��@�S�ɶ-�,��$�B�[-��!����/Riن�o�p��0d!>��"%�o��/&a�ۚ��{h~�4��XO(~�
'�A�*Hم�|ݐ�)?z�p���ΊO)�q�MN ��2Dd��C;&�F����D��1���@�v���II�����~8�f����O|���q1�Ms��J�Ӣ�$	%k���9f�B��)�7
y1��wЙ*=�E����SP�`���\#9�A���I�� ������?bݦ���wTY�BJP�Z�}�S��ڱ�F�a҅�[G�y�@�i���*��W��]�(���n�ڇ�d��fX�*�\��*V+mpS�k��?˅c>��/���Q�_�Ԟ���d�G���1���	����'�q!���n�.������(l|�d[�c�ԗ[�UC��s��l�y������B���⼃M�y�so*�H[L$��{N2/4��ezoܭн/�v�2�5F^�2�F?IZG�!G�k,�A���NN)�gU㓉����&��P��Ex;�%H��O�b��R��](����2}_N}�f����Z
��?k���r#�'J�e�Ȑ3�z:߳��3���o��;:,P��B]�7q\
5���������a�u 'Iu��f�o֫�"�	Y��=Xz������
��Q�7�z�&��Y�m鷭�Ӷ���w�)OU�R��5���N�5������C�>ӴN{�j9���[��k��@�m
��E��P|������Fw묑T��=B�`ۢ�c���s�>���!Hi��md��|��]�F��<�x�{\B��W�>$�x(�8��aV�A-(j_̠)g3m)��E�l1i(��H\#��"�B'ٜ�Zr�`Ltp��%6��[���V�ɞ\a�� �2I5�؍J���H;~,9�w:iP��٢�= ���;�	G�U��=p
�u>��Cko��oT8�J�pp
�iS�]W��sS�#�07��m�-u�C0Dv8:�Y��U��ȶw8
Ƶ��0�G���Y�4TD�ǅJ*�����4����m9��*I��>?�%�Ƣ�\��qH������Iس��PNc����$��[!���%#�4��*G�k��5���@,[�5����֒��G)s�;\�s	.z�rR��)�Z/狂.׵�ؖ��ma,p�\*G7��%=z���@Q%��,��3T��� �b�9g닢��>�w0�)����t�oj8�G���;��6)M�{��q��T�L��l �8�﵁�R���F���U	#��;Ϻ?�4��]h��d72��"�`!���+�]���W*E����Xӎ����	]f�� .~�Cً�ZN��ӗ�ݰ��Fa~�F@
�b��ϔO�%���[�����J��j�ʢ�����c�ј�����E��$|JN}�PȀHJt��#��@�XcH5¯���u�i�̠f��H��� ɇ��CMc�m���&���j"�b��ڨ�5�%�8�R�'�:�mBcZ�L����#�����j[p�����2��0���\��ŵ"2Q�p�����*�kn�^��N	� u�䮥϶u)�Ů�G{)AD���lS��?��mJ�c�NI�ڡ����aq.�:�x�`ezO,�/XV}��rFe��o^�������3������	~ة�ԇ�ӕ�cަQ�"��ށV�M�V���#{�h�W�R��qf����~�=y��F��0��?������	�5K^9Mt�a�B,�M0JO��5�(m�qG�_\���i��yh��~�q@G]��<%�	�">ɱl`��׶�v֚Kb�)B�NO�^��b�'�o}ԙ҂��;���'C�����݃��Z<"D*�����i{�!��s̽�&i~$�B2.�Mf,v��!W��	��Vg�jh�U��nR���"�s���{7�~̸\@�"����N��P5~߹|��5~`?�e<��Þ���ܺ\�r4?�A�� ���z.��T�Ć��vu_��:�s��o�����?Zqg�-ܙQnol���k����>�II=����Ƥ2�C_y�߹]yzav)i��kTq�w�G,i�&tw�+k6��!����]�*�n��go���àZ�\�~,�̚�;�]U�,4����a��6��m�@֖l��a��:�ԕt�5*��ޒ┷Z�l��V{G��s����#�r
���	3���wB�?2}*#�$6.���z�50D��0��޳^��,�˭~C��y���HPvl(���$DXk�TU�P�)�w���m'3c���h&����ݤ�����p	�$G����T�o'4����D�!�=���6�$��v���Z��A���5q�U��6�ñ��?U{.��e�T��
Ӥ�f��N[�)�}U �X�)���n�#j�b�^����S�q>v�^uI`J���1�c} ?��"�s�oF��h�˪A��d�9Vmdnj�	8a��,N̑������$Jd�5���q��2w� �RV|���EVbQ�8r�M��. ��F��^���鰆^Ԅp�c3��u ��V1�EWVֱ�=
2=�Y9>r��/r���wS�ɑ`6ŖE��G
�H8�g��*�$*��<2q�m2?`<]ߏDa�Bzj)6��=/�i}�Ϭz�Ŗ	�͇\h���
PZ�7sR�kh��? ������3�R܎�p�yn�>�-�ے
��F��f�����Ϣ�eiw��t;\v�==�p��T4�0iUcz�(�8�\�/�1��eቄ���Y}�e�ii1=�̆��B�V��+�=y��ϛ�5� ��sF���vϑ�Y+�V�QZQ)�IB�=T�	^_�C�(U����6�3�m!�{�`c/��2�hɭ�q	H������|���epL��
nV:�7,f�II�k 8O��#��? F�J[5S�-ZeF��f�O ����=>݈*>�%#uq��^�5���׽�������<}�_O��h���F���]�W�Ѭ�w��뒟����W��Y��b�#o��u�d.NV>~lo��;?T��Mj_	�7pg�P,^�2lm8�
tj���S���+��ڟ�M1T�Wx� �]P��"5yC�Z��.C=� %���@�қ�mD�"�c���vo��V2���-�"�$J=�{!�Ȣ���{)UG�/e�7붏�0�U�8hoT)�(���!ަ�uz^w[�ɨ�u:����3�HT��3)gDA��}8c�m������YDP`1����&0�R1����|;�HX`�M'F$b$3	�zA���5��!�y�T�����<c�W��W��Y�e$\����V��?�RS��۱�E�+��gUd��ƅ�>J(�W&KG��5��Y�D3�؟�E���ĸ�9��frn]��T[��]���� P��zݯ�_���:ҽ{[ �3���g<+a0L�e	�J��̇�E�`�]���I��4�a�g�럎G�J�BL��Jq�l�|��A�$���p$�z��=A�[袣�&��H!��e0�Z�ٵ =�ɵ�QEc��0 GS�Lی�<�<���'o� h�z�a���v[��<� ��E�����BN
���Mu�Q&�Ԏ�0f�W���/��V$���� �C��fI�����un���#���{�o�
�Ќ�7��R��u���G ��۱pL�ڇ}���Od�Q}a�POa!nzu��u���sf+�����Ӄ6��i�A׎���N�0�p��΍����"ȷp�S��V�e+�x؟�%��gӹ]m�D�	�6�t�b��I5p����b4��r���J�m��N��=�}.����c�!s���i���xȦ�Ċj��e�DK�Y�zD�~�2�FJ�ӟ9�}{��v2�@e�����;�E���e���=����ƀ|�RqTØi�SJӻ��
۬Ee�{FN�_z����!�P��`jޝn�sk��hW*|w�)�(�٥��(�L�z�s��ǰ�R�	�i������G\��rw�1�M�u����a�����`�+������xx�ܖ< �)�Z��(�R����:�#��2�����8�4} P��+fM{������ܽ{U���)�~??�/@Ǡ ����~P�*	�.�$DO��c/ �v&EH����D�m;�/NW2J)�[(�nЕ���﩮$zNI۞O��{�vV)v�ӹ�Ց�7��;W�Z~��b+}�h~�ȝ;-ˤg/���/�I G�������?�N�VG�gJ䯾�]]��+1��q�R��qf�WW�*q���7���R<�K.�$^.���Y� �c����{n�G�$��5��s��6�7Z�ƛ�cu9�wC�A� Mr��)Q�D��R���#|��J�#泸kG�J����˄J_�'�@. �y�丛���YT�Xp9��o
9�����j/�L7��v��/5�ބ&i�r�6{�1\��56�~G(��(da�?�d��u�B��Ŀ8���;Z��x|��ؼ�".��i�����R�%C�p�ҍ���?���oh/��O/���h�n�8 � ����2%L�b�j' �х�u� �L�W:���B��F�o��V��}@�k��b<Wx<�{U�Ч&ׄH������n�Z�	��it���ɞ-�uV������ĸ?�s1��l�;�@�H2�!9�ľ��������n���k稾&�XU��n��3���J쎙['�'�k�)�^����B�Ԙ�[��A��Rk;��\W���au�;\��65@;�[G�� ��>���;q�H�\9�u�����5�h9g}�����=/� ^����p]�Ss�,*��'+�*x8�')|���-��/ZS[�x��T��jC
��FM�[��ҝf��1z��GfS���(8�<�Zt�d&W>�f�@l�bH4��v2���Jy��Ū5��Y�Rr���  y�,qs݈�`��|)9��ʛxɍ�"G�d�˷�l����#,:$�Ӯ��d)X?L;,� �-�fn�����˶1��tJ7��CP�dP1���-��Fm�w\1���04�� .��E=���g�g�E�gE���B��U Kq�������99�{$��aᐔ��Nh��
���"kTM�ެ��e$�c�Q��F�(ȏ�;��6�Y�����%?p�%�(��
����MG�@uiT.���5��ⴟ;og(*�p�A{d��JF
�_"ݷ�)M7�76�x�{���_�*���b��v)����J�B��3'��#��mB�\)��	�A�v�p:��=A��㓱1���)�8�����A�ާ��k�n-�œ���]��/1uD��<wI�Ι�MTE�ȼ��<���4�5���Ɓ��t����m�\���j)~��D�ZR���E����`g��z�|*9�!�!�>6rpTwE~�%����Q]����c��V5.�Up:맺eRa�7ҋ=P�ޛR\C+$�!�5�Vy��@�fŔ�k��EN�M���Uc�����vYI\$�)@Q�����6���9�;5�����&.�.���.j)��n�N�`�)�Щ~�m��{�,-)�7��eY({A�q4����Eh@���y@�e~��̜O��fWJa�]c߼�t�����h����S�g*x&�Hp���W5|*�$?��5[A�?��4�ҕD�,����^�Ȑ��zt7d̡Q˓���$��s���=��A�~��Dy�eCԣ�C��[^]��]�d��+e}�-���,����6��F>�厠�S5����t�"�9�g�=������(F�(�j�Wh܏Uu����F`2��F����8#����v!�b�G������d �*�\Et�/b�X�o�;�is��#�5[1j@�V��j�홷2E�J&{O�	W�r�fI�
�*iɪ:5�VV|�9�ʰ�}'�IyE&g�O8 �=PI^�@Mf�c���#�'I��sݦ�m.v�ľ�Q>Dw��Hp��R���ڶx-�ua�F�6�
]ʟ��:��P*@YuvQe��o�%�'����	̹nx���B�_b�)Sk6%S�C��늟gmz��'U�5��!	�T��2��������:�L�W��� �����#�Y�(��@,|j��%��M�!O���a�Z�h���khӅ��H{�lع�DE�?q�в���i$��u���U����͖��MU�X_J�I`����̂Hpv�����BmjAA�+����m��;@���_/�{�׶Y��ȝz�52N�7=4��ظ���\<����`�a���b�O���iH'�o`�^M����)���g��\�ݝ�����b��n�?�DvH˭�6��ЏIi�4ն`�g;�L��p�t�x�A�!F��숲i;�(n<��'����J�
�Ov�o%E�L�O^�=[
+�(*��V�~��$�Wih}�t����?��9�f$���]��`�߂1%�ⱌ���EZ+� ��1RB�T��6;�+,z�aU�M�G=x��9N���k��U}Q9q?���qX]��F�m
�X�db�[����]ZÖĘ=QB��)�A���~����3-�[y�0����u=L#bs֡��B$cܔ�F�]�/� =&��!Q�W�y>�Y�� EQ��c����r������)�s�픎�m�+�R�7�����~7���-mٴv�,���� �J���� �*���&t���ߟղ?0�mMH�!?��q@Q'u�L�0:�+ƥ�v\�YڳSm����8�Q�F �4G Ngl.��pӕ&�Df�ڪZ�r)/I�-wĭ 9vBu�	��<�?�e��<^qC���Ү�1�n>9�j�C���orpm��o�7�E�]mp�z	p,����t�i�&:�ʲ�h���r㣟]���8��Z��,��
�
�'_�1
�:��=�U׮N��%|cڞ�Fn�Q)�_�kB9a_ �|N�z�����G�SX�2�h�*�V@S�jG��k����|��(Q�d�ī��ҦWl�E�?�O��g��áI�Q��� k�u�g�D�E��9!���"��(���.�!oee���4��D�0����]gj:m�L�='~��(!���vq<�ju-+��%p9xfa�OՄC�3���x Q�C�l�l46P�o��ȷ�u8�:���p]�ܓI�/���<X�|9���2wl	���AT��a������'��Q�I�D�V�%ϱ_e��TL���e�,�Q2۴o�4����y|n�d�'f���j^w��8fP\�5������
Щe����?v�#�O���#g��eo1�[_�6���_:���N��<�~�w{��Q�l8���B�����5o�T���f.�j��L�`���P�3�mu�����R����f��;{���v�c�G����r[�Nיi�cu���Zl��T(^ �M9�4J�9��>�Dg�����ǔ:�%m7������'����
�-�N�����0���;�~��0�,�H]F�-
�Eu7i�'��K��{��p���9��X��]A��n�"�;��uU�Z�F_-�k�,���\��/q�f��ړ��K�_�q��w��c�_�D���PPH�z��&���p����U��մnyAt�+�@�z\]�K�Nwe��D�zX�����pEue�qI*f����7�0߃����<T咉Z�٘�Wv�f�$Օ��9�z�Oh��t��3ۙa+hr�Ũ�3�OW���hR��[;���^zi�O�8��l�����K&3�y���x�Z�������T&�"Q:��
iEJ���V>�ԭ�(��8����VnC���%M�����E��GSǥWj��U#�Ig�^�b�%�B�aHz~5/7=~���h�����,C�"�U��kD��ǒ�k!� EZ����"b.Q�aVgh�؞
�4 3O��I�fyֱн�A�ճr�LCS��5a�Ȧ-Xq��C��Ec*i�%�0o�(��z�>�BZ�;�;����7�w���B�{�+���C�>LJ�̤!�(_��&�5��P�Y���Ș�7rv�|���$���޸_,�^����Sn�m��u0!Ȼ]bT���l+_0�^xX�-�0V�[���q�E���T����'�d�^�}��+lYQ�4$
�]{�
�� #JB���v-y��A�����/l0�S���V=	|�ŉP�F��U6�����`�W����^�z3�XVz���^������`�Z�������sa��j�3�L8�jᛘq�74*p>���B��t���������s�01GRou���'I���~}q <�%�;*�fG� ���D�<�cQ~��)p�m�n��m��	�m�l�IتW0Dw�z�2a|G�𴞭Ÿ��20e�\��<��dA2G"�.sn��uhFg��K�A�s{�Z�%�b�?c�"U�Wi��n��$E��V^�����C%4�~-m"�y��&�;�T������IO6q/kdkb �>��1���T�F@�sP�Rr��v���p*5'D�U�p�z�	0Tta��y��^�}�.o�DM��l��P�T�	ȃ@�]���IG�\�!H�X�Ha�M�1�����;Q�o=�''��?�Vp���ą'V��9�t�1hN�$?JkLhG$}w�I4�nM⮛1>Xo� ;(���-qG���=��W5Bq��A?�]�J�|����3m � :�Ҫ�K�1�ܵGto>�gǙZ�˱@~�Փ�t�&z�Á���-ςI�~'[�9n�N�8D���0�"�:K��2������޷a��mK��[���XT�_専�!���i����_�l]#�#�&,�/Vd�ޱ�X�܇(�%�̾��'���ʏnX+"��s�ï��h��K������/��2�}�0@��%mf´V�̎�&�*R�_�j������8�s���Y�{�n�+8�*5.M��Ki8>��z��$s�7���HG��7�.�F���%5��'��~��	e�2ڈo���ޟ�k��Jgo�_�H�q�1ڋj��y�c!pI���q��ǂyd�l�1�X6�-����i�֖):�Q��AW�WS8����s�r������/,|kR��P��x�֗*y�^q����1����D�(��[Y�&�i	�!�s�)�r˴��C�4-�Zunj��Q����Ib���e}�v�~`� �lkO8�~�Z'?ˤ�Ɲ�T�7˫��]0��c� r���f���ݒJ��Kv�\��%#�"�o���
s+l�R~�,��Ő�7x7�<�"`jӟ�O���E�$S�l��,3�7P������k:�;>��;�#�1��k]�c���&!tj�TA��>|�ե4u��/��7	��)�fV]�.��w!�<opV�0�K��^�\���� z�h��_r����p��za����GH[s�l=O�ڿ�ga4pW�����Ö6��Wq*���"�=5�&APJ���.�D��q��7��-�D%������b�3p�tl�]������v.�)���?�?e�H'G�k?1�X+MAsux�2I��4 ���9q�ԔR�1+5b@�n��(�>�_䙵��_P1/@�M`I�s��P��It0���;G�\`$)D~C��x<������l� Q��ˎ�,Rآ@��s�W��4�=��(j����o����h�+4�E�7/[�y�[h���=E�K�ǌV�8q�r���k�tr���#p��ΗF��0`��W�L�q@�q��cvL<��F�A=�)��-�i�Z��{���+p�;?�Y��xJ�Il�D#��h��	��c0�h�P��4���]��*-�O�۷��c��� ��Qga���a���Y	<)����\����Â��Y���/���ѧ�9sZ�/H�c �Eٟ��پ�:��Vf�W-�@�״���\���
B\e�(bm��%�ӱD�cb�Y?.�,$[,�W�ZÈ��
�J$�&
xG��A;���_We[Α��~��Y���c�p
K�������3�6����ɒ@~C�\�+�U��B�[f`����Ѝ'��Lj�`L&ڞ+����s��>�ĝ-�����СuiL3�c=���R+L3o��s��^������8��`:�	��i�(��U�4�G}�����J�!�h9OHO( V���k�C���K�6��:���п��Q�^s L>?�!����2ޕp�����X��R�e9�rM�>����!����Z.er.��a<A��;n���cB���&j�P�Ʉ�W��=܆?E�/G<��"%G�8}|��:7���������-�O�dN�X�5�_������F᳢{[t|-,���q�ʔγ	J���>>ga0p:�����A`\:�Z[{�s�G6�^g�i>lQ<��9�'�������I����J��I�:tI{Բ�K�za�W+h����s������R��|\q�_W��p	���~��8WQՒ��}�f�x}�g8�*�����1Bj-����N/Ȫ��):#�B$����.�>6���O%O��jL;s6�O��9W;��i�����`+��|m�UZpڭ�/���n�"i������}k�9�f9�ΜY\(������fU`� ؄r����K�|�����w'�'fM��@_z���7�']�T�&��WK�͂�e@�'�6�2i�$�Ct�.M�} ?ZĨ�nj�X��g�/Du6���|����5�$�ߧ"���GͅB���.-BG~�[��@M8H��Y�̖�;����'[n���C<���>��Eq�b����Q�Ch�hޒ�p�
L!*�M8�E=n���g{R1����!Z�z.��=1*ps�<��I����~L�EB�g�+��Mr'Z#ͽ]�q�ʻh,ƞ��myf�	�wS�[�㼵�]�*,�.x�񦎟^��y�xz���9C�M�� �:�?�� }���<���ωC��)�X*�ܚ)�����O	�3��i�_5��?p#Y����U���Q��)�NT���1�nQy�*�S��]�k6�J�luI��r�Pte����{<N���$Sf�T��Cq�
TrT,�����¼�z�i;ں�w=yY�7�����"�zF�nTh�(����2�sIP5�
6��a�4�E0>��q u�p�c\���L���v9ޖ���="�^Po��%���]�2A\*�!fÆm9$S|*�&E�UWz|�et �S,��ǚ'��Mᬼ��^��JR�)���ө۸�BZٜĳ�J���M���eN��H�ä�� �xPJ�1q����Բ�`��?��܂�dJ�õ��'@S�D'P��|��ub�t$�����Y3�L����?X����p��?aW%��߈*���g�/E�Bd_[�&�~yK���	����n�}���UL\���2�G؀����_��Z%
{W�/��.�����~����g�B��e�:O^�t�q=i���L��4w�������뽞��X(��̼>8�e�]�q�Y�ֻ���Hʙ�y��������S@��uR��IUc���X0q�YU��}���A�T�e����l>�vIC���q0(�6�WOS6�@/�v��ĸ8��no���	�y�����:�Ȇ5!��5 o0�N�~�{k>w�C���!<��5���"�[�Y�D}�ؠ�Ek
ܐ@���I�V�å�6�jpd�MQx5Mg�Ag����Ⱥ��q��[��$��T���&iO���X�w]XL#��T".E�[N_f�\�vl�%ھ���e�S��q�*E�����>u�4K���6N�%��iӛ���L�z7���2��\	�cN��z�u�Z8�TyL��##�j"6��;����lcӇ9���������E��k ���z+�|-��p�Mb5�f=Ο���ߺp����^�@���Su��#�aR�42����\\��ݫ��أ?� ��B�y ��a ��0N�����D��=��O{si-{\��$7�.���S.>��Jcc�w��3���+$�ɗ���KXMp�-5@ē���{[�K;a�+�ڀ,��������ㄙ $��eI��ډ�}C)�䴓o�o��R���#�C�5�(ƞ�{-+���N��Ɖd�03��U�T�J[��Л&���o�껌��3�jƧ�nd�BM�%E��G�Z�`H�������� ��.�ukb��>����Z�v�@�w<���~EjA�1Ȗ�)~��ޮ�fDb���t�.�]�ՔR��ɹ��4&�YRs5l"�y~��& PK��Kۨ���^#��b5�$A��S�b�~7[�����j鮓m"}$����ș^F� �[�տY`��S�4�N�c�v?�߆W�|o��;j��t�����Lu���JտFx�q�^����+�
���=6��"�䈖��23K[OwT6��mx��+�����}ȑ>^���Z��J7�A�)�j����RۙO���3�|�vi���D�|a����.b�+��gn.\����Ƭ�Qa;��N5�«��I�#��D�v�b>AI4@BFϊ�����3���&��*5,M�]�\}P���@foVJRs���i�ߎ\�
��yK��RŌ�I��mZ}�vJ�	+��Ų�0��Ow�x_�8�@���}��N��A���A���ݕ�"ƙT�<<_�2��L4�&�w��~���� y] N�H�J?\p��_ȇ1a<[���E��W�JعiV)��3�-�@���fBĬ���.�b/3عxz�&�0	H��Κt�b�]��&q��(�/��@��3Q3��"M�����[���h��l�%=�����M�PR�$���A �q�K׭ЀRQ�;��f/5m����Ћ@�{�n=�GI�2;a-��N?@Q�v+�^b��~�A��v1��+}P�G]��x0\��&���J%w�#azKƩ5`h�߭�s/^f����~�&O��0=L�)ҵS�O�WL���%-�cY܈V�U6�#�`/���%l�%h���A����;�cS�U�u����@-��Ϩ<R�K鍟<�%}���GE�|�RZj��x�QuZ�u����k���դP��]�
�Uh�:�T��O������༗�2�-��7a�<{Ue��2��� ���d�5
�6�܈@_��e�/�o��lA"J��^B��Ve�h�6nW#��\���_�� �[`f���#V�7��yKi໕!���_,k��D�x���B�����{��r�1Cpi�W=���k������zi-
=�����K�Z++�}�x��n�W̴<7 �h���M(�M�s^��_�S���'����W���4��a�TQ�����{lc��"�T;0cvL���T��ed5�u��x�ԏ%WG2�HȳJ�C~��{]}������?��N�u��6lN&OZl^�P�vI���D�DZ�M���F�����\�DΣ���;M�o��9�P5�V��Ć�|����N���"é>SUPY�&�Msm٦
{f�����:�}�.������Gk{��R"A��2��^�0t�<p
9/�E��X��}��yh��{�K�[�|*� ����hTGJ�����lQ���;g�I���y��%R�۬|˧U��bRW�k\��Z\4%m�V���%���S=�Z�~\��L@����Ƨ�ac,�]�h͵����H��VG���,�:�{��mQ�D�VG�x��WFS��2 �(��_�����S�t�=>K�[ �z�^Gv���g�R�vg��R����@�W�j���<cS$Q����9�h�?4#MIG7�{�f_,[b���! �a�L���;�w��1+K�F�hnz�X�W�x���D4��=��~�Mz�4 �w�ʗ�~���k�n4o	dj_�)�����{�m��=A��f=~�ٕFT%M��$�X��^O������k
�CjvH�h)?Q��Y����l�z}s1�}��&���u,T��s�c5ys�Ջ��׻���P�|\h�I���j���Y��QA{:\$�6����N��(sv��3���ӕ��>��Y��F��N����*�6�o��S�����ǂ�wwl��I���5�;7�� �_�f�N�m����ف�e�~j??��s�Ŷ�'S&V�or�@$�a�9�9�>X(���1P�I���^$D�/Ơѿ��[k0���n߽k���S9z��6��p�����=	�|<"���a?o;Q	st.�� ]�|�sP�yc�3�����G(�MaD���Q�TaJ���ޖ�w�X�C��/DR�*!φy����y,=__�r_X��F�)L �	i����4�r�
���
IdO�N��.��Cٺ�������I%AVd�UY�7,7D�]�1ܧ�H����P�NV�E�mj�b��J���fZG�sl�O	/���{��"=͞/r���w���4��g]�F7���l�����5T���2���V��51�L8N���>`���<
��l���y�sڜ�����҉�0 aw��m��,����X�yD�O��i���qeV����W�Y��0)v{OG�>�u�nvZ�S�{�,-�o���O�,}u!��ui7��A��{J����CmX��+-�h"m�,�,v.�����e�U�r�*�1_}�Ü����.�ڀ�zs�V�k�E��9U�y�����L@�-�8%��.ۤ�x�R�6L�AV��($��+C*󀧃~֍'�
�ޞ_���|:��u���@����&�U��T%�D��SRt�#����s�:�m���'�K���?X�ld�fg��s�" ���*ɠs�Y��,�wd-�	c�[��!���'�T<�-�$z�9A��!����� G���[�	Q+��|ɡ�0BR��Z�,��5��g��`�@|~��^aA��5"��b�Ӣ>]������� cG�:1�O����Eb�}E
�
���h�p*�ŀ1�ͧq#:�!�YY�+��P���^�ז��r8҄���4� ��r�@�LCS3U6���v���ҿb-&A�C�S��4KQT=4�&��a�r�9������6��O�+�:��LA�UI�i�e���24��rc���e�**�!�]1�NL��O�I&�i#;���S�����������u�u���K��C,I�M\~&n���M��\�^����p��*~�x�s�#�Ӷ�ua����s|WY��޵��xŤ	�R� q���z������U3|E��q���F��>�#p�A����j+�V�=�R�/�e"���('$\�s���&� B_ʚ>�2�])�	K4�-��ujWO��*Ѧ�2����q:^��m���t�B�j�pu��H�� `���h4����ŏ��~h���?�6����'�fNw�+��rdkɭ�a���~�E��UhB&`� x`�Z�&sa��R(��p���xHS�<�8P�^[����K��g���W6&\�Ӽv���7��� �^8�[W�d=�Q���B�4�[��0�lK^�N�.a�DZ��I�؀Fi=��IY������\B���O�E�h:�3ЕoL����c�L���(B����I��AT�y�#�S;�@Cҳ��C��B�ջ�1* ź�V�����j�Y���O�����=���Š�@�\����%�ޅP��&�lMt�߄�t��Ey�0("Tt�#ڪ�ڍi@�wਖ਼��)��l0H;!T�� j,����(�o5U�������66x�Uu�Dz�?L�N��G��ih����lWx�6d��I���9�_�qB_�}���F(��d��R����#��zx�!˴�h�I\�(X>�?�;��'J��l1l����wd��Z��y��)ͪ���2����4k�H�b��j�ݝ9�
�JY-�cn�Av�)D\?0���)�#����|����L���Q&�7w�[����i��aƹ�b,dzp�������qJ�-ې��s1�I��A���&�Vdń�g��_@Mi�3�f&�4`��o�RȎe��2�Z�d�)���|=�B]W!o�I�,7F��d�L̺�Am�ui�b鰕Q��'+��&w�ϷR���b�!G�Q]�=1�z���A��~�`��%����6-����qM7�g@�;(�?�[���{�8��cɋMa��DY�8zRp~^�T2���&mm��P%,R�bO���&�5`�����F��a�t����a�BbpL��=19�AA��g�	���L94��/�D�nx1(/�?�����]���j�h3�q�		����t��a�7N?*}��⩵�S@g��q��mup�v-���a�L�,�i�dW�W�+#��C��/���`d�<���}�y~�M�0�z^5�E�4;�8�I��9���i2{3S����{UH����1g�@��)|�`��Wip��SX÷K��c�[�\f� ���*�D���ﰦ��iѣ]��;�yX�ӿ��ܙ~!���}{�7jag�*ʀ�ПW�>�C��d-m��&G܇�K�����MU�/�Yש�L�O��R.�K�;�G&��.�(�mxA'�pg��y�i�9�1u�]�N��M�Q�q�7�Bh�0�HRL�Yہ���GK����57k���`��S~P)5����"�p����Zeƍ�Jɻ�~���#c��U6�@&}�8�y#j�WBC���{�ƫ�<�M�HxM8�1�-U���r(\=��s�K�Q.3RO�VN�5��R���o+�3/�L�dlB!5d�zOL��1��V�!�8��К��%�31c����.|�Π����9�0����(�

~t�2=�QR�BOKJ�W*"雷�@��H9�"&��.����z3)ug�U׭�>Q�t;~d��1�Z���E���W�T<��h\=<��ic�$6�&�V����t�(�G�t�{Zc�]V-�At������i�zLg �۵h�&+XPL�:X�tdKn}<��c�7�B�{ŕKq���"�l�H���4HIs���WS��P~r�"�R��+�Y�TqB�G-�g`[i,b�C]�P�E�L��Nf��ޙ3�J2��/�5��2>՜ݲ���!f	�V_`�Yynf�U���QI=�x0d���r�@ˁ+Á�H�b�����}J�Z=
9R�*3>�ȟ��6ZE���]��)D���w��6'H��4��<��9��ܒ�Mѵh�²��`	�����_��D�JN%��g[W�+����Y,{�%�5����V�Oa��,�����\���*�/4m"v���B�"]]��]L
��!��訥��s�;��������kf̨�6�v����(^���]j>'s_�Y��Zq�Z ��;�k3�N!@$�YzP��H�*����1r�+�Z��eYf�+��=&"�(��{��U�Zf���?�����X��#.T�um�^���)Â�-�L>�G@"�̼N�Ϭ���1DK�n�3#H=�"0j`@�OțV��U�;�f�#��G�5�j텴ф�]
��i!�Z�V�;��R��xdZE�� ���%db)��v��Nv�O>�V�qͿ�.p_z=~S:�+Y�j�~�7x��T=�GY�7�h�h�,g�q�ba
*E��^#��V��H��m�W|ְh�]�ڬ��D醗c,��"H�jl0aS���?���w�U3�?��7�~wA�ǣz�9�9���цCE�|-W����汆v��6������ڗ���_^�g�V�3���$3Bg�e��6�d���_w~x]���(��S�����i8�{�����z/�Ȼ�Z�#S5m��v����j�/v�����Vb�L|"'h�l���]����U����?D:��@��lkr����ݫ��7��cْ��¡e�֡���({���[�]76}12's�U��ܫ�����z��c��,ŵ����!���^��C��������{%5�d�>:�z�_�
�����*Ҥʷ+%�8�*�mE��uu�z��`�X�;�����Y�a�%�S�)ԻN�mZB�4�
h�Ԁm��Qf���b8ӿ����(Ɔ.�u�4�Y�T
�_��BkM�,�d��-�`"#�GG��T��!2�S��=.x p&�="4��Lf��p*N2:�����\x�Y�~4C���t�O�h�G������Q�}����9F`�bߍ�I�����ov�Ǘ%9��!�6�XwjL�䘱�7��>�Œp�ޱ�;ӈ�U�xnَF��Q~ѻ�/t���tq�c���$zŤ���}��. 	���`��qĵ��^��x� (��n����vJ�4,�N�M�U�"�M���2��#�GOk}�~�|xq�n�����[Ĩ�ǽ�]To��B'(��{��?>�Fix��_S{]F��F����O��əa4B�n�D�x�'k�B�rH��<S{�|���C���?�l���[!ޘ�x�m�"
�5�vJ���^��7�����CF�P�Uo���=����um���yd|�O��	�<��P�떠�8,c�	�-g$/O1��g�ob�/�7c�S��9�F�L�a��e�Z|Ëz8��:��5Gu�yJ��MX݂�!�䳎���{�'z�0�N<rmuxJ�vܼh�����/&��U�/��x�����p��1��2`��l�/Lg
���-�gY�� �ռ�+�y����U���ӧ���Sch^UAu�\0/���H.��KŨ#s+����A��:���yUf�ӿ�biz���������˵#򖴣��p9��� �g��G�aOvܾChIa=��2j�����?x�4��
D��M�D1�E/�%����d�3��p�%ɴh�LpN��x�"�fr�ͅ���\�;s��hR�X�^NI����U�4"!�SHyaN����>j���]Q-ңh��F,X擦@��O�2_��i�Yy=	��!�����ؿQ��a$��}�s���j�l��O��6��"J37�ߴZ�#���5�"��[��֤�#����l=�g;�B{�w)t�IU�{�m�T�8;�[�FJ���@�Ѹ)���&�S}��2��Ȟ<�%�ϫ[�B[�+���o�W�0��� �w�\9��
=�-��"���׆Y��e(��n)�(����|&G\�n���F�c���Q���As�]��7a#��@d/Ϛi3��ٝ�GO���F02+>c���A�+����G�귵5�>���i��+��C"�ǥ�B��:Cu80��w�5�m!��[���� �n�W|�����\4���Ȗ�֞�$����g�*�����*^�����;*��]���]�ӭ8I����ے��t�L8����qD@Fı�F���h�#����i�UG���P�_�����ȿv1�]�Y.X�Z,6{�4��j���|p �8��Pe�s�Υ{�X�l�SH�UgEMߢ@E��8�7���my�J1�>9f^7��dG�w!�]V� ES�+���֥kXSa���g%�9����"@RJ�$aH)o5�40�w0�G.�`ן�Hg"��?~zㆽ2e�Q�����ʾ#Vm u*U;htr�	�^}H4�0
�
�]Ϫ�Ͼ��w�2�Sx�E��2φ5,��L�4��¶y��i��9�&K$+��L���J����H��ǫ�,�z��d?W���;-X���l�[Vߥ��h#Ib���N~e��Z/%�c����o�>�>2UD�B���c���kg��e�H�K Ǽ���L��>D�^I�Ew�
�(�+.�6�d^�Z�:k���`ޚ���[��)�TsbN�)���ͥ�W�Lʳ�Wt����ma X^���F��GN���`�:t�);�1�r�}O��CO�6���=Lc���8ƥb|:-]���f�-C*`���cJ��;����&i��T��s	(����10�qjr�{ O��q�1��]���6�p-���o����sǯ�6S�����)L<��Tt>��4�F��F �\�p�)�SAh�����i�18��C4��ҕcSU���l
9���Hk.X1,�A�3�m_�V�C2ޏ�nb
ͽ�u��U�a����ɓ5��u	�h1�'��g�|Y�c>I�����&�an6�� �5�E��D7����J�ϖ��j
Z䗨Ӑ��%�ٳ�@�m�{O��!e)-#�c]4[��Z&1*�:�(*�2э.]�{pU�`�uU�Hr���-���_��u�5��.邮�6�R��i,&&�
�e}٤N�]qfk���Þ�������,��w��pA*���$M֯@�N?�T	�ǊB����A������x]���X8���G��_оԎ�'�+!r���pm����_,��W��Cf]��9T��VmSe�k��L���Q������ҎּY6��I��A�қۆ1}w�;5�n)� �z�8�0h�'��-�Z�u5}���߬y�z��iC0�q�g1��]Ci{Fm�9�ӡ���H=lj���a��������l�b�`�,�����ѣ��]�ɉ7 �����k�.���ʰ6s�~���ZV�=[y����z�Eo�T��4"R���{+*���r�0�r3[8�;U�V��zV72#�Y��� �"%QZ���ɯ.�5���g��U-0�B��rw����:�(�O5f㶐!�e��f��;� ���T���ľw\q��!��� I��(:�H1|���uɋdď����p��j^2,\������gA��}���4�H��+Ff�����s����+x�>��#����򀘨�3)��q��7\<X|������m�;�;|�pԇ՜�4嬄��v�{#�H�*t���]^�N VP������a	�J6ޠ��	\�
N~�p4Sm7��&�A��wx��c����-9���*N�1^Qx-rsQ�kec=�$�𗼿B��P%�T�<Q�ܻN�gu�;+����И�?��3����P�\�滇-RI��*L�i�}X"�' ?�=�wr#�)�ϣ�Z��أ��2p�B=����{*.��c�̳�A�`��:{��-NG&�7S���d�)��89^�y\�)���:�D�eM��V1�.�Qr�d���U�G���	n-*�j�Tk��Iv��?���*}�9�\K~
�*u�P������1����g~s#ez�Ii��X=���=�I.9BDdz�M#�в^#W��e�ӀFi���JA���KR�T�P����X����׿(�J,��d!(L�C7J�n��Sz�ar��n��'X�n��/ןu�e�8L�O��O��,�o�E#+�M����I�cҰ���@p8�v胪q�簆q��!.�RJ�`e({,}ザÞD[�4��^��� �9ác�JsKA7���_��%07�t��|-��	���
�65�2�Y�6�w�Vj)����G<d2^�&>@ �c)3��Hw�eUE� +p��ҥ�Z��C�埱	Ҝ��#�C��G:�( Q�S��|�#�XV���Xu1��o�B4zr��%�8��CtW����\�f|���j�܉����Dn����SqX��q��T�3�ni亣I���re�� 9#�̒���Y��r�_��K��l�q����f��;hZ��X�A�[l�#]õ��W `�B5�
\�a����6�G�̱?ir$P�@�6��,���]@�š�Q��/|�$�Z`��%7Ϳ�n�2b�<O����������k.��>#���q��O�@�Y>7a�в�=��v�/Ki��y'g�j»�O*�H�L�R��;��q�@�~f��ז��0�Ƃ���d_�9��$ N�3�NG��-���fy�ެG�L��Y���{tT���(�\�O	==��^�Y�7�㣡���2��tHQ|��r�,�����������/gb�!�_�9�?}xei?Fi�SqN-��č�CY��*�:�j2$zr��� p���*�n4�@J�ύ�I:בz�����'�`���B^bL�Z�pI/4�����5��I��Q�Zb���7i�8�,l��^�Bhss2�4Ȍ7:���\�{X�����($�jN��0��5�[��l勘���0�	|f�`q�?��$M��k��g����Ԧ
��2C����-I���mH�ұ�P�י�l�|�;R"$;`��=eG$+}Č9SX� �E��%��1�g�TG,䳆�1m���o�@��X:�,8@kLD�C�Pc�hz-��K�C}���#��
}�z�e2^
�����
r�=��������%H���yӸH��k�@cY� (5�P<��ҽr����W������U���1Z����KC|ߓ���2i��[�81(/�%�v�G�>�q�d�8H��B�	w7��&��OeÆ�ۡ�
b�14�K��c�ʊ�5�L�M\b��2�bx�$q�,�P��*SqNd�e���
�[("�lB"���$*7�^����1����{�/�D�&B�{�����]��!\�e:0�}��ʢ�pD:t�m[��8�Δ��
��yM�'@�@N�����駠��MvS��U�ݠ�>�8��H7��W�k$U���4`9��!W�{wd���5#@�B��a>	N�#Ձ� �+��K���ͼhCY׬�hy���ݰ3���C�T�l�=)ޑ�LbE����X�}Nd�J�z�����>��V���yRI��^ك���Ā<�ˢ$DԒORf���D��r\�*�g%(�wrS\O�}�%�Tt�����<َ$F4�R���M����m\������(W��QO9�Ӓ�
I2<��^3G 1�)�3x��Ud�]~ ����Lɚ̡���*��8�]�z�V����8 [՝�Z$ŧ���f�AXNe�@a�*޾��Փ79gKHK�ݖf���@p�D*Ls>�5�g2���=�Z��A4`�ǧ؄㘬Br�3����F&l;nO�P���,ի�b�PQ�ˠ"Zv�{��R6�wj�7DqC#CԵ�|��ʑ��Q�Ai�*��J�P)�H�r*܄BIZ��>�hǟ�,������O,1�f�e6τu�](;@jn��1����-?�D F�؟��ă
��� G�$M�[�)� �xa�{Ȭ8�t	#��k|�&��Q�� a�݅�6���S-�`�U`�e9Uw�93]^�Lݕ�DTɜ<�F��c�^�8�j�Ϡo����|�vol���
�$�Q�� Ϣ��mC���V�ܠ|������07�~D�>�,���
���~-������>��	�*�{ ����"d�D�����8���m�b�;��e>��Ӏ�4dukMzK��TLc����D8��U��x2uۂ��e�!�&�>��w�F�*6꬜�w��!��"񦐄޶��ߟ1v&�-��W87oƙLo�=pm���	zn��j�N��Zy�ص��"��E�ti��P��gu�#+�� .c�쓭2V�J�}�D�oV�Zd�x��-9|m��;�e���h�$J;2�,����J���~��<��[�e0h�@{�b�ծ�L�2��d��yp�l��F��Vב��N�0������p�C������n Ԑ��PzS�:���B�8��Ժ��x�>+��HM�����I��	�E1bO��]<z��2
���\�DM-!Ĵϗ5%��w-تјo���S�:T��3���,��+��g��D6+�#+��s�}�Yx)�q�\�9- [Բ@[P!9P��c� i5B�?�
��K8n�o���gT�����jh�>.spe�q��᱓t����ȃh`��>B< §/�_Nȭ�GzH�� ����)���c~����Fn+k�T�Q��j�s��V������[����>��i�H��`G?l���{ ,�"�f��C�Cཟ kN�� ��J�ow�`��/��Et�5�� H�6&Et��#]��V��YȀ|a}ㅓ����'�3���ōPš%ٳ�#�P^��R��@_�a��8m$�sA�Z<B�-���m<TDnԐ_|�@p��`��� r���.�;��VK!��g�ʀ=���4��R����oV!��f�),���V��h�n�EgJV��Lf���PaX������C�w��5L�I�n��;�7���ֲ�����nÊpu�,֘z{M�ċTrVG��]1�=�b�R��H'�"[vl���x�_w/��M��ژ�+���֣���c�4��6���
�+�/��?��l%���&Pa��H�"��(! l�U��Ӻ�Ms�JÜ��q��$��� ���=�I1:]�/�{�:�ਖ਼�<^���2��.�_�K�yR���7��D��������f��\j�;��0�e��T���6@���ȑ�"�ucbB�}fGڀ ���rda�7F��Ccb�]ۙ9o��Q��`�d�)������j�� ���s�C��q���Qj\ՏC���V��팢�q�X�P�~Y�`����ƊP���vN
�}(�Gn\E�����.��v&ow�A�`�����^�&�E�ےId�El6���)N�S��D@��T�*-�����-���P���B�36���,Ä��/��؉��`�p�<T:�H�;E=�2�0�ȜJU:��yǮSe��(5%p�=����-���*��E���X�B�x�b\�}G����A�M��&tme����SYg!��b`2R:pʎt�X��2E&'K����>�5X�nX�� ����+���9d$Ъ��w���i+��hR�cCC?�*q�n]̼
cg�k��,�<YFd�hh=Hk���Y׿H��Ң����=|n&OĐ��2{P�ȡ�
Z�&�"�4�(�[�r�q=�'���;�ӧ�?�]��Aeq��Fy������쳑���KRU����"b��%��y�]�U i������Z��H��}yT/�����,7�v��ZJ�_5�m<N=��	��baN�*���4d�NG�>_��`ôީҠHb�`�֜v;�W_ǛM��-{�藬��)��*F�<8��z\��߮)��(�Է���7�7�.��h:�5��XӔ���+��
��3��a��hå
�������`��PA��o+��_F��۟Xᾶ3m��-ol������������>�>���E4F��C���}k������H���N��1v��j�j������1x &B���i��p*�+�:G���!�����/*g�����j���WM7Q�]�r�4�� r�O���HR/��,���i����M���}��`�;[	k�<�?^�צ
�9�����]L1+<��oi��N��b�{-�d_t��k��%�;�9��P$��.�bc0�w�j�幩�"4[���F^�1Ji�u���Q�Z�g�R���\�p�F~0�@�u,v���>L��o'W�-OP ^��wN��Q)����$����p����䯸 �6�G���w��0�k{�l�n�i�(uY3�`e��	��U�u�vM�.ʹ��^���p���aP|�$��T0R�D,���zE[el3�G ����y�.��%�XYKG'@�4��c-������z�'_\�)Z<9�\w>k� f�[^;�v=g��C�!Z�����|?р��	�m�F�N3�-׆:�n�s!��
hq���yk�A!)�^*Wl��vS�q.���W)�t�F���C�Y�"^��Z6�js�ub�%nʻH�@7,`��9]^��_� �a��JA��W��;��N-=��󵰾	���3W�rr,�yon�@�LXo�1�_#���;S�![�sfv�R�4;�t��17��Z���7��9��4��]�R�p>�BO�+w���4�ZK�.6��*|%���m}` ��I)0��nP���W�,(�������n��pACX�#�'��oA����$S0�	^�ۧim��m��^5�9�tVg�ѧ *�e췑J��f��vZn'���+���@s�4�G,	����"�z9��{��&<��]��L{����G�g�$���8��<�*�9�����P��I�i��]Γ�Qo��p�|��l��-�ח�>wr�O�շ�yy�����\|]�?WM���P�>�M�rC2�ND�	D�/��&TD~�;��_�_4G*��rz�o�T�I��_I���%'z[�Ry���u,m��ĝ�t �%h.WDUj��3�;�IV� �_�l~8�OB�ٷ0����v�V��)X�R����4��=�7��k��Nq�k�LaЏlC빦��.����������ҰD��^����.��^�OK=�,�r���4v��8�4 ]�<OE��j�WV2��ڨ�֛��-i{�Y�l�ąȢ�jo38�JCN�C�<��nP��3�u��O���O�V�q!�p�.��Ҩ�)1Q����UJ�AE
�Q�f'A���e�c�,4�&_���>6%~&ݩ�]�U��l��V���
�:k8�'���Mr���P	�^�c 8�v;[��������P���ZҾ��u n��S����6W0�'G�6���t�b����Z�^�������6Fy����ÐI��ʙ��F{��*My��Ş��?z�D8G����>.�Mw��^�aKi��*��Jy�n��y����Q��K��� G�a�j���XI pr��`t�g�a���L�ĕ�S�UY����m,?�MaaEr�����A�z�5T�lI��\3��5�lG�ƛ�A�п{���9��s{?�2έ,9
�``�m�:%�=5���-�E d|Jl�(���Nj̾?�k��v����Pn�@�S*}��sE�1ΤJ�l��|��J�(rY��RI�v���؟�8���{�^����t�_�++�u><¶s�,���Ar�q٥�8���ef�`�]��>&�0��1M_�U�c�l�u�G��M�R��������CǮ�f�Z��ϫy��ql^�~�����kJ^'�K����8i%*�z0>��L��_��7+w]h��%c�\��������P���AGW{��� �9�hid�9�r �ՏyQ��o����Ŋ|��^Yc[�����$b������h��Z��K�w.��mnAG¢�࣬�dZP��#ViBR5������W��D��5�+*c�v3ACK�-:IO����3b%N9�>7ځ1�;�O`�?UsmV���!�>��3|�[�Y��c��lf	�'�P|!�L>���'q�-P��Q$%�o��l��4{׏�a��f��?NZ5%�j���N�,�o�[���b�e�u�6X��ra.�V��
�Jd�����\�$�?����6Ĕ���Y��#j����8x	5�����eO�S�.?�����m@��]ޅg=��$;�H����K^��q9��1J�ԟ�{��	5�D�@�-r���#7j&�rq5�G[t������>� �����㫰�l�ѲE�="����i�����6w29w��>���ATATزJ2Jbt):Z�Ļ��u)+t��W�u�ѥ�R�w�d����ϝ�ȁ	���}Ӌr;��>{�Ϩ�
לUR:5��!|�����)�7��`t��+p	�
&S������4K�԰1��`���J��S�c���$������pV,Ξ��ݦ�!8���&��ڊ�e*\�(�T�"�|�[�6i�tܲ�؄U&~��ۣX!(�X8nE�qɠ����v�����Q�W�����n��G����b�X"���՟ݕ��򞊴�W��/î6B��2Ӯ
d��AaЗy����+��s�֖|Ff�}�Qy�"�ZTE�q�e{b �¶��0B�S#��msV�s�����W+�
�F�v��hw�E����46e��洨歉���ZR�@|����<\��Ug���'b�】aI-/��9���e����ysRu�x�l�);�}Q0�&�\��zɋk������>��zd�`�^	�?�V��`�A�ܫ�wCơ��#%�c������T�)j�5]����
\���@)�B��:��(�J��my81�1n�J	:�����:x��0��68�ڙ���%em��N<κ��_ޞ��~�ѱ&�TcdW���=�
�7�1 �/)>"���:V3��#>����#"�l��$���Q/'j��"s1r)@�C*��O����0����h��/M 1v��ZE~�`��	`vè��7zNV�k�U�ן�=uڻ{pqȏ�(9�'���l��l�=#������]s@ɽ3U,�t��E:���g��d���<g-sT�r�;Y\�u��wV;���7\
�@TaJ�E虣��0����6��>p�.��xN�P����̯��=�7'u�\�y��! �HS�+�t[�J'��Ut�9dK���sv�+�B�[�5��N��F��RE��6����!�H�}@�g�� ��4�^�Dq֘8���P��m�#��wx��,������ �T	�5N��e�O/+�/��WUt�sƷR\� x<���LE^��K�\��0�Dv���~pL7,ʭԣ��!}E	�X&�F~���e��_�b��L��!������@CV
Kz2������;��vV��̥�޺M�:�w���-��
�4^�=HV%��^�� b�8m��x1-����+�������,�9�N�QI�����7�s���y�m2Vb���s�r_��,��)�D��8�J�C��:�I
���㻶%s�A����ʸ���G�^��#�����%.}�m�I����۰�G��[�o�?�Bnv���;�F�l��p)Q��D������9� )�t�MUB|+ _<��۟�$�hi�r4dEI��u�eքW5���v.�
��ZY�p_��Y��ǅ+L%�5N�ea���b��2 �AYt?x���	:P�·('\LW�cS�㞮��� �5b,j����^z`g!��W1o�)��9!�c�B�L��6c�P!�T�����ǟ���@�/���n��H^�ݬ�0a."�k@��Օ�|��/��`Rrd��@N������l�V:��bt��-�_����Z��*\�.�~)T��ʶ�B%��5�P�q1���jP(�b��Vͬ:a0�aيҔ}Æ�b	�����P�h�'CIv���s�뵶�Ҟ3�oNH�%W�h9�3Z��:�
�2�̏���P}Q��ѹ���R|'q�������a�]�5�b�!�.N�G��Qa(���1�N����@C< קּ�P����%";�}߈-�gK�V��%����t�������_�֠�7b ����}��ɢp��N?��'�����B�,!�a��G7qW��ɁW�����m_��,+Ta�C��\Fϲ#/H� eNz&�3@��4&TM8�����>WV����^�Aj�A��~���w���X̫K���'����eƽ�k ������_6hJ�/J��6�@byHYK4�����F��drw�����Qn,� d(`�-3DV�(��o�9�E�d����8��l�F:y�|�[HU���u�wP��#[����3�3��W��{u���G�e�a<[Ŧ^�
�MY�N3�Kp�Y� k�[V��.[5�.�_Y#�)cHA��`�-���ON�)һ��\a��k�_)U.�u�)�c�b���/w�����8��5��	�D[�ĥ�+�p��r���K셠Pt����>h��"�{���d��>o�  Z���?����)�j0Tv�|��~0�W�m�RS�K������
�_�:�/H�����L�}�P�QD���,�l�&Ŏ�������)�С�-���S��5nvc�S�|g{�Q � �6$H��P��2� �[<���mG3k��[]���4����
v��ZW"�C�Z����)9�!ép_����d,>�� ��>�Q:�| 	_�]	&Ô�!|-Zv�3�Ҕ=p�\�j��b���.R>�>��3�/ۢ�E�V$%�v�v����	�M���F�$$I�Y�c�'��92k��$I2�{v28��W
�%1����W�t���T�I�^�s�`�zܢ���r}�D� ��接I��a�+�|��We�e���AH�ϼӼ��y�3x�i���(�m������xqP!�/�|�m���<�pot
�a��������SBr!��
Ҽ��򀮶|���k#lD��3�O�
�l]T�}���D������u0��0n���3�޼}H��@�eF��2�Ȍ���B?O������^���s'�J�����D��,���_ ��ޫ�h7O���ўt����vU"�]���t�N�Tf��1v�Yɦӧ9�ũ�n< ��Y�<���X��tb�ǿ����q�?O�d������r���}i��O����a��+�C��3�'6���,�hb�S`p��F��p|0����<�������ʽ;Y`��P����D��ZaZ-&}.뢻�ţ�e"=m�:�3}�BbP7�J}�U��M�\��J���:Ĭ�#2|f�D�A���$)SiVt��By�ɟq��L��k}�h�n��j�V����펌j�+�?�"˥Y�Ǿ��1_�@��/H�[�*�ڸ+�$��<G�A�SBic�JL���N�����w�!�s
1	@)�Ì�c�3��^������Uq�$�kիak�ؕ��P�p.��Zh�D��j%�[a��@L�N�m%�0fH����N0D2Sџ>�w��1^±g(����vday{�(V�n�n�P�V��M64L��- �%\�x;�MI%�u�ҍ��>�E@V�-�]�ֻ�Z��!���=P��F
a�9&���pW�@|h�k�dLY���n`<�7N�Q�"tvF��-Tn��� ��%���;'_�(;g���W�ڗ��[�-(F{f��s���&>eC���a��U�w8 �J�ոZ DF��pP�f?�$_B�0`��K��r:���2�>� }�r��xo=	WG�����#����M�ա	��t�	֙.�L��LN�vh[M�Y暕����(Fex0��Zj��"`{�n�	�̦�B�6����<ͽ���$#����0YWUI��R]�����c�p�1�<BnjO6�B�+���������c���M�|�wKG_}���Ǵ~ ��ܷ\�J��-�pj��DN��d���>jq��kՙ�VS _�9���Њ���Mɥ:�W��*�
2��Y�		�]f����Fk�:_ħ2qS�шy��2ꨣd���o�%��Z�,�t0%�"�hx�X�T�'=��,r��������RS��u�M���l�x�B��c��Op�?ds>�>:�;ִ�ȓ��E���;:qHz�;9U�h�*Ô�l�]�Z�gX.$��H�D'o?�w�J�����N����Y�!C����	8�n�;�D�J
��ӌsu +��J��&�V��4�CK�}�?��z��<:W�'����W�.�?���F��n��?ՔR�߃'$<��ق=�Tvi����u�����$�%s�-����(��BV3�W��?���p4�FFy'Z�Vw�T (lN�Dp����E��9A,l��
�V(��K�9��t�V��2P�C���Ĭ�������T۰���i���؟�M��*�~˟�ݳ��o��+a��(�db��EZ؍b{J�*;�4C=����Ʀu���Es%7���{"'�Θm�:Zd��YB�R4[��@�"D���d�Qz��Mͪ�T�h�lś��
3	����T�K��c4��f�O�?W{F����m���fّ�:K�AȪ�����:��c�q%��v�_V�=���Q�����gh��4������Jϓ����ǎ�l�arw q����6-����z�< ��O��n�lx�|�9D����	��Z�[-W���w����/��rh��%�l�kh�|�As! s��������&��A�r��������C³⸸%
��W/b��7��+=�
E�\lTlF��|�p��(�:����h]H]Id���>��o![rq������}N���%����|�� ��_ǭd'�Ｙ@�j}�oVۋ�jo�~�r�yʍ熁7�oFe%*X��F�ޛo�Bw�9��o�&m��v���(x7ťZ���4YțQ����w1���@ϳ�x�%����Gs+�~,z��J�;��v�8T���m�1KR�]��xF1���ā"�ݻ�F���Q��������H=��@h{������_M_0�p�܊J�[��m��95� M)FO���HZ~��eBS���4b��/E{��q����	|4J�~8�[cp� ��ө�,�-ۊ���^�(���+��<?��_
�V�f���B�K�ք�ID"��4���pGr@����8��s T��[�v߈=xw���zd�
[���`��e����p� Ӡ������(
��{�;9�aW���0�.�\?n!�������7��|��oL� �
���+ͣ�Γ��Sw?$�����6T�p�!_�_D�T��W�;��7�7�,W���XX�޴):~��X$s'�?��gI(#8++�J��8K�"[������"�zE��h�b�)�t��	J�|�*!�zYC�(�z���YU������DZhnj�/��s��*��Y���!��M�Z�s5�
d��	��ľL"=��,aĚ�����|���H��qx`�&e��j�1�qKq���n*��+ �'�5�^�=���g��K���°��}�gf\�`rVЦ�����V2R�,�1�����BH��:����hE*s�7�	�Ԛ�����u�*S����w���r3�~����K�G(W���u�z<K�1mY�Q�6�}d�Q�kgI�2��J�9��.��,w��jlo�o����9����㘦VD���2��a̔������N_)s�ˑ�	��(����.�Q��ݤ閡|�0'��e���)d>�6@��A|a�ו��[��K�ǃ�`d�C,������w��z%rw X��$͗��7~�ͬ+Xğ��#eJ����9Q�6����&un���:�)���zۮ�	?��F�D��b&m{ϢM�H~ �G�UG�� �~K6�˟Gj]j�Me�`��i�lyS����=	Ih���1ˁ���w_�#�Ǯ[ݭu�A�guӧ��_w���O8�R|с�@1"i���&�mum���v��?�.!cڧ���4�toQ�an<����u �4�$����{���ػ�n�\�PQX��daa�֢U��7['2�Nݧvͬ��0+�������VQD�K�R�/O@����8z3$!'��g�g��؃01�#1�W"5�ٽ.-S�z���K���K��������-�e��Kzq�@b�&��	����k��Dʻ�xy�7$���Ddl�1����"�B��_�H�>o-��g������B;��}�a�S �#��+P3�T'ֶU���7�<��C-+�$bJt �JA?��_���ȋ�?�����2_tz�����^�?��d�W�Q�����Q�m����ʣ���z�*X��)���~�Ð�F)��=�����g�Id�_��\A�l�p�3��i�Ɛԏ�z���[U��/�l��^���>���Ț�u���1�a���%������#?v�"��h��e*}/�f��ү��l/$�*W�m�?�������W�	A�7�n��>C��^Lm'�s���%nU�%O�5�@'�;�E\Θ���AOeFu"��я��m�%PPM{�6�N�:�Aǘ�<���$0(^��Vz�0{�Ӏx$S���	�/� �:Q6�qwTpH����;%��
�X���?�]/�}'	V����Ε���gnV%Ov����s����m�"��^x�}��[ip{�u�Ϸ�>Y�)��a`�-C��T�K&��@q���$�`b�lJ�C��Ûq��P"(v���܍�N ػ��S�szv�v��p���t03G"��Q�]̵|�Z̢����k�˝�R[	��h��p*��'}�od���l�`��[j� �*�rf@��n��������m�Z7���u,�9���ۢ�ЪN���M�|W�]�Q��1��6����c�A"g������.�&)2� ��9�dm�g8:� �/�}���R���v��6Dê8�0��k̕�}�a�!Q��d��+�\H'��T������s?:���6� 4w�Y�z�� ���D��\���F�,�[���[��/�Cզ�L��S��*�q:>O�\�/u��8P4ȡ"D@�zqz�>o��*�Jv"��Ӊ���Z���<�w�si�*!�b��Şs��4�ͨ���cR���~�S��bm�MT�[b�ȋ�<���<�����k�V��2��M����[����^
m���|B�çt�Gm}��$���/2��Ei�C�W�:�R�o��-���L`�k�E�wh��8�������ǽc޸�0mU�&5����5�;��h:(.��_:mǵX	eԋK�99X50�^�K���oDH�[�HO��mBYߥ��x޲Q�BⰡٰ4��~�UtJ�Y]-iX�D+B5�Vc��7��˘��C���F60'4ZY�zt)��H�.�羰��oO�gFuX�G��8ߢ�`:��N�zS�;?�}�ڰ�=+4-Œa����#�{/����,���;�@�)�������?�%��E&���&%뽎�J���S�.B���? �"zj\-��#:~��/%~R�$N�涅g�B��&�l��A%��5�S��X0�W�E������{$rn#N�������Pl��̵����%L��-��^TA��[��+�-�^���O=�ߏi��#>���J�@M:ݾ�/��r*y��\��V�xO���*�|~s��?�0��^Em��ZeiX�AC *�0����\V��� tg���;�G�<����h������XV<������Vu�ik�E(�UAL+����Z��uR�v3
,3����ځbb#��S�`�\�n#�1��3���~sm�dg'e<=%�F�H�Ʊɡf�y��	H�͊�Q �y��Ƀ9a��k��?��^�r�Pu�us�^�����
�dlW�PQ{K�Ԝ��ɭ�ɂ��nru`�p˨$��\�^�����K�A���7�A�Wk(�!}��)O�C���1?r4_TŬO�J5J�e��7E�����^��yƨG	|���\ulH\`��{��8c�`��r�:R/�-)a����WIAJ�/�{�3C�;:��y��>�Zj�����ڶ�ܰo����?f�
��5�����С�R��BWi3O��T��yu��դ˘��"zR���֭�dz��6K���r���$x�BL�Q�4y��fۍ��ͳ��Z�r޾��pFv���I�t���_�0�ߒ��fu��ƿ��b�F�?�)s���XD��м��啌�j�?AG@	�L�)����&T�zY�1��sst �J?�p"{m�`�|U=�ܭ�N夵��b�h0WNTi���e9�l��9X��|:H�?�W���p/��D5�����*f_��N������C@W�p�v�v���2)�~�:��-�`���F�'ю��E�]�(�A'���ƥqp�*i!���0?��*���O��_��|XZB��ɓ��k�I�A��j��הWc�&���G��a���z����R��!7�:Qu��ܜL�������P�_B\-��ay���r顣��������h�RP�H�S�H�g83,��3-v�����Q��E�)|#=�3'N�b�5��Q9!��4�F1�Gy��5�>زF 3�3$~����Z?Ҭ��(ʠ�ݗ# hN��$%.=��Ty�b�)��q��MY���(�7��H;��[D�������(T
 d�: �a`�x�,"U���!�i��eP=�T�`,���04T�"�n�'��E�����A����4�?��X����3�Խ�`�J���8y����T`�kAu�������I��A{8� &��u2��N�(�͐�a��u�;��S_ ��C����9�4�����݇2D^��YS�?4o���Ǫ�$?�=����H;\z�}oF����"eQ�\����Kj](C���Դ���\Ґ.``��#R�(z�]%��YL]4��?�4e�����D.�3�-R��&�<�1�N�Z ���f^i�C���|��ME�r�B���C�nq��D�/�� !����bqY� �Mz��9\�p�j�k+Yw�]-����h\��S��{{�X�W���0��ѝUtq.��^���?�c>��� 
M�'޼�ߋ#۔�a|������A>�P��Ԡ-�Q�qa�gu�ao�.lS$��}
��)��o�̰)"��v��r�΀�-"�����H	�{}kgh���K�-�'�<9i��S܀���FbXl>����H*����[M}V	������K�����U>g��\9^����.S~��,7(��sa��n�#��Y?��@*k]��P+Kn����~���<��3�j�w�^��-�����Z�d��F�7��?fZR��&V8��׸��	&>`� ?�@[��lNV�N7��D?��V����q��O����:�X���LB�W?FM]��f��I���M�Z]�m��cٖ^�9h��{�_�򯥼��d̶�h`h�#�Ч������iF��iGy,�ˁ��P"���$�=4�?D0lDn^F���# v���p1@�	a];P�ɨ/	d|>�.�vC?���s[P�2�c�@k�����^�A~��I��MtݠF���D�!�ߘ�ɽ%�<�^(�#�η�X��SC�I=0��X���D⡧���@�+�>*�̙�'K8��(����x��ߠ�tw�S wϔ�
m<�M�MN����k|z�}$"�t�Q�<2��	��]���G�_%쁮
�� �7���W7�8 ���{����w%Y���͹Za���<2��x-58�8k�Q|��Ǆ�7'���\�;veWc�*�,��2z+:��J𕫫�z���{a*�m�gltB��f��)I��G 5��[����gK�aT��	�]����N12���I�j�h�q��`�u��Io�P�՛���sN���o��ϐ+��e��*[
6��߹�~h�m�z� �/��ٖ?��}G���Ŭft�8X"˕���N4����r_�ݒ��k�W��JFb�w���**#no�$}��h>X�k�eS�G��1�Kc�.�ɓq�o!7�յ:-g&N0�A���@A|1mJ��[����ר��s�g�V�O������{m�F�x,�82���3��������ݘЀWÇ��l8M3g�cA����ۑu���X=R�DC5�����{b��rc.�w�\�

'�KF�ū($A���(X�0H��{D�<߿=��>oL�e�\��[Fg��A܏d�L���y�0É}#��6�~���hi��t�.��
I�5tr ��a�<(�i�/X���pu'�9�sb��g?�_-��;�e�dVcJ{m�6�uV�=�%���L�鸊~ ;�,��a�Z��x�W��� Y�gF-�3��,�#*��Mr��g�I���<����\���*'
�ĭ��ߡq2����������Sk3�	D:V�����ޅ �zd&9��O�Ԥ�^Kn۽B�a����	ׅ�� -�$q�-I!u+�[̞3����_����"Bb.���RT��B��8�F#�d�\����ۗ�*���D��H]/����ϙ�́*����i� 7�55\泘�B���&���h|TC��U�9��#M�=K���A̢�����_k@/�)��aM
F�3�p'�k�$�2�c
���p�
g9M#	��W�E�7Z��$i|�^�c�᥷�|��wQ��Qj�h▀�%�t��Py�w �Ő{���0�d=W��j�*Ȥ Mk�����^� ��$��uJd��:�R҂��r�苭�����N�x{���&�!�l����l����EIG��p%�r��8���ƾ��P��ד�F��ϼ.N):}��A��1C��OO�~�����٘��\.kSa#Z5~"�ФO�_'mޏE
�vڼE�)'`T!��:_i �$UXC��Y(�0���3I@t��J���	�Tﲵv�g'����Q�|	ʣf�X��Eʉ�?�V�gq��uL�c&($iN�:�WI��p�/�8�J���������E	q��IJ��?>&K�Bż�# E;�J}������R���O�=�n�;?Q�d�O�% �Яo�V��j��(BJ ˑ�9sٙ��݅����H��^+M�GsO�R,���?2$�\�8��̄W_R>yt���� ڜ�F#S2]�C�)EZ�p�M�m8�N (�Iƻ�S¾8�UC��S���R�^�٣��q�f�$����#�QW8c}JB!�g^�_��_n�(��%f�U���"��S�Rr3�Mz�X|b���b�=/��Qn��F�^��z�})ԥkd Y���Q���)Yӌa���Ruy�)XO�i��?���#�F������Èp�:_ry�i���������som�{�*kDë$o���AV��jsRHe���%��X�׽��n��q'M�Z��ְb�y9��7��M%���s�:R�����z*���� h�m}����ҿ!��ڎ}!X�}��}���2�ӹŹS�ÐQ�\"�d�Z])M��F�N�NѠh&������Z��e��U�t��8�#�tb#���1p�VN��ߗ�<�V2����3��^�Ӝ��6�]��n�'�����	c�{cu~�&<�^{��	�oh�^]��:Z��RU!_���۟�sיw�g�g��g���Q3_���������ו=���4����I���Uw��Σ��H�>��n6g�(��苶�p$�'�y�U��C=P��[�ӖO0xgHvL�ᛷߟ<��E]�C"N=��Cs��즱����3�n�Wg��1�9�谉9�t9�H8o� 5����ӡE��	(��O�Ff�B�e۷t�K�=�98�.�������Ԓ|6�#rX�:�����.�rP��E�JD���r���0���-%+}����@�Y�o��I�śWt���꼸֌�>9Q���ڡ@�q�=9j����Z7�v{C��}��]�G�ܦ��Z���������w�������Aú��BO?Y}}���K��o)�d���Lfs������[3�vw5�П ��
\"����A��ڪl���m�{�)H��S]���7�H���8�F�;��U'n���?-$	�ix� it�t$��'8?ԧ�de���(�!G�"R���Q��7/�[�{���Y�0�W����� 6���:��a�L�\8 �[�k�QOf�y�@��5��4᱘����N�2`X[�R����������y&srwi��n���e+W���`�b��v��@��@��w�������N��$mh^�s����u�e�S/�	ՒqK�Y
4Y�]��j���N�&E0�B�;���ڛG�sg�C+����W}�N��K"߫~S�	�RJb���c�G���
�/@�̆R�}ee*�� �.�1��b�<�T"|�� �T6�y�^�#"]����w,��L��E�����15]Ŋ
�M��d�a��,�)ũFqFR��%w��=���m�T���zٝ���]�_��P�ò�>	��GOa;����5uj
�Jc����:��\��5$\���ӊ�D ��F���ks_f��5zb
$k#�lC�zJ<��9C���Θ��pa��η����*�\�8�p�G���MN|����v��IQ:6mP�f�[�SFe#9.�x\�7��r�mV4ᱥ �<ﹳ�f/��)��؊s������j�YɈ��!C����{iI�kEj2q��k��Aa�ǣoT�� ��ur��pE@���$�2�"3K]%DҪb*��:��۳5 ��M�<���9�Şs!�L�U(��a%�h��K}z��4��Hu0�=�c�!dk�G��F��CG�*}j-G�nM�s�98���΍yU!��, ����d�g��joE�5���z��8�۫��0��IA���z x܇'��*�����d����T`�ް�h�`���[�H�"�Q�M���B��嗢�%��K"�*+�n�=~	�I��j�3�|�nm�'*�]*$!2��[�8�m0Q�U{�@ �d�� RD��Joiꉖ]�=�kt��:�7헢���o^�G�O�A�a�)e��W�.�hY��t�'�`�v��d�h4@囤�F��z���A�8���MĒT��OP��*m����U�~ocT2��(蚧�Yo�`r�Բ2�ɧ%�1�3%��S���f���X����`tm�Y,��Zy;����U�/4��z�ߞNw�&B
�;��D"E9NJ�ίu���s��Q��f��f���Do������{���|g���s�m����=�+���H΄��z��G�2с��J��6���=\��{m]�HkσrH��^�ɤ�ܘ\���H⏬)/[��9��c5�Y�7�X1q	W�.�D����	V6�\,��|���X3�<��*�3��}(k�*�0](��(Ur�!\��5T�8�Vh�D!a�.�Y�n����3��U�K�Ya��^M��h_-�����p�0/�m���6y+m�����p�a��)� C��!x>����&rTh4�!��0eP1$�g�$_`<^�ˑDf�.�&c��8��~nE5>���y}�R`i�r���^��V]�a�#�}씀c��Y��×4�\yxew�J�U��Q����F��d���b:*9�ڴx�gx�s��M�N�6��K`��֥`晽���@؞GdJ"vJAq��Г≐�W4 E^�ݔ(�R�&���:jM�X��k"���[u}�l�!�U 	E()���@.�Cl��J���N6N#�?��WDnzv+�r/�~�}�m�� ��Q~<��I���ojn,6���ٷjid�B$�D���c��`>����g���.*��ZѸ�F���/!�L���;��Z�h@"����iϧ��a�O���"�l'x�/:f�"�����Y����&#"Й��d�M���ħ;כw�NT�}KAm�ްJ�&�������)/Uas�Q��/�X���&��~�D��6�LZ'&�H/!g�ϟ!Nڅ�����$��I3W�R��H�*MR���x](}6�(^��_e*LZ��[���g���&^��L A���4$���~ͧKt�f{ \���M� 0�8��Ĩ�W�d�nU�W'�eu�a�����1�f�8�}ʪ܄Dz?#�]d�\��˧��!��S��ufm���Y~��1S�
I��"cD�Ǥ<b��豒��$w��`�ѹq�zI����GBU�~�q��T�i�w�,�dr�L6�H'ܨ3�pWv(��u�O!f$o��ӭ1A�m���Lّ<t���.�l�̆l�-oP�C�8���h#��2���]��z4EW=p���a��_M��P3�+��R,����>6�����1K��t�Ǌ^�F��2����1���}>�1�6x-�$��Um�W��I�Y'G,�����5_�r%�J�ѷ���Y^<��� �4��'m�"==Q�0�w�>L�kyW�x.Z��r.+�xyV5��$]	�I�����RF�3��%h9��}� $Pk:q��_�)�e��'U�#!$��c��)��x��a�#?&6KS.SK���[ �ɮ��W�&4��4����3xY	����:�g=_TV��a��YT�=���i��=zze����L�|$:��������I��|E�:|�Ec�:�D�`#Jm��ٳDM�'�mu�x*���""��E��)���\@	`��t�x����U'��}��j�7�|�XMvַT\K��6<�(�L
�.��_
�@���h�Re'��k�/���"a���t&,JD~g��J��4ڴ&����Ms*TP�p�Yr���
*�:�_��V��7R�t����5�~���o�������=�F�oR �O��\dK�|�!�t�m���s��ഈ(I���	�� V�#*��3[������O`W�ߜn���Ԝn[���rv�QC�0���u��چ�T�)�˞I=]B�p��$�4h��fP��ðxK���'/:óe��PeV�hk�~��m�;��8@承��y��VS�q|	�9aZ���f�|�D�Cj�����%-��Ј��$y(p�/�h�)��O�[ǩ亗�ގ��\M�MG����yd�kz.N 0ԏ�݆���?|�L�'��:��~ő#���X㿓B8��!��z�Jʛ��t��}������t�6���$�+�����ɟ�m���)$Ufl��útŠ�35��GZ���7܇��1���g���n�U����`�P�AKYĽ_$����Z<�ȏ�	<^C�坒��+�@^:����j�]������b�q�apRpO���Z�%dԗ�[��"�ۛ��x�
����9����U5ӝv������mf���o��F��iW�xk�G�M+���)@�R��2�R�u��x;����:��w�h���:��q2;t��)��]|��)O	uK̢��*�ۏї 	?a3l:>jxK�8P32[��*(��'��6;CN3�~�?
���ua�����綶��b
�2��B`
���sDrLQ#|����s�;/�Y�sW	�X	}��5� �=��9(=WٸT��#�k���l#��R�*�c��>���J�&�ݏ�~-n�~$t������U��I���Đu-�KKm ?�j=՞@U��	�%�D�,V8:�����-G���Vy��Z��٪8Gh�cͫB@ ץ�������?���w��Oj5۷�t�	h���4U�2>�_�����p�5�A�?`�R�K��86p����Z�4_ߐԺ�z@��'I�Gq�l�X��Y��	�)�y:ޔ���[v�^p57�O�h�zh�oAW�a��P�`�����m^����7�b}�@E��A�<\�گ���ߣ9g���~p+t�<~D#o���1EN�g/�V���_ez�-�q�3�@��oX���ؙ��:�a����o�`��fi�����J��m'Z�
����;0��G%Ք� FCMw���{O�qF �~��Nn�-¬���Q{��kY����c�,��|����nlg!j�{+	����1������ P+6 �.��b$pإ)䭻8qu��:�\�H�Y�v$�ة#�~��jf�:�F${��w�e~s��w�e�Ȃ��k���sɈ���Yٵ ��6M��&A�E)U�5t�TS��\�w<�#6�@K��>�
fi�H�8��b��6Km �<���Q:z���sK�J���Lih}���p�l��5@*�T7f� 3�f�vE�����~��h0���NK�������b'8�(��>�oCӐ�M$�∞C�?b56�Q�&�����x	�h�O�UZ[#È!S������~ oB�D��^���dD�PU�z����Q���/Ug����<E�"�gL�\*~�{\� %�k,��׈� D��+��e< E��t LN9��@�����o��LyW~��!����h\�%P�h����f��}�(+�Ka�3R9����Ⱥl�(���-��q8�8���)C�\��D��H��7��}��"�M�ݵ�jS��j�(�Y5���B:q�I�̓�aM�yN9FQ��˛f�!_��u���H~8?IW��� ����@S�ca4d�P�\;���;+��V ���rAW��¯�>�ړi��ʁKj2�^^hY�b�N����H3
�<.�Y���x7�zy�(�����7�i�7H�߬��k,���is*��\�{�wI�lL2a;����$P@��FD�W'nք���|(��Le�%�����U��'y[��M����cq3�#CeS�[��uH2sM�□�]+*�N�9��F[@�%�)2R�dFù�>���C�'X���� _ w����A�zC����Aw��mΔ3�X!u|�=�W��q�_���q���!�ewB��q�B~��)�X�McXN��)�"����(�8���Q̡�:��|Ov��N�/r���j,����^Fڣ�.Y�� �m�|�ݫb^O���9�>�����9m��L-�H^����g����w
�5�bͪA�^z4p�@�.�zb6,+ӎ�Wg���������D�1h'ʖ΄�?FN��{��R�_&�d;�t��UQb���"������r�H����$_�q4��Ő{2�X����qT��t��ح���c��܇�&�b�Ɉp�Eo��y�Y[k�U�t���Ӭ��k]�]Dhzlbj�m����n�?_u�eq%��3qZ~�[�M(G�u��f�!�mU���V�n����*�'����	o��U����Q�2㤱��|Ym����C�s}m��O~��\�_L��tV�=;H�Co��;�n��98s�^2�pu��E��X�Iê��D)�up���ВؑD�`�uL���j�7E�WQ7��Q2	i�>̻��Mj�\wh_�?�YmeTH#���}����g��	�aJq	��A�J٬�Xܱ|�4��2��$�rhc��Q��HU�9?��0���Q,�-���!P�fj¾�.w��%@ޮ4�_��f?+40���V/�c�EM�aa������`H���5�?�tUG%���Wo�j�FI8Ɛ�g������Q��З�돸��,ce�s���9��=?�����3[%��-͕�vE-�*�g��b��-A޼t=T�Tc���O}|$[��w@�
uc7�~�P1طR�3���[�Ū�i���Kc�1k�r9.��*WM?��ǐ��U�P���Ƥ�\>f������z4���o�S��7�5�{�m{҄o�!�+��B�>��Q�n������e���*e
��DĸXH�zg�E��Ө�t2߱rG�5�[J��oiNUb|Y���/�Ө3@Vne�w͢uL�E�%X���yr��GqC_B�C��]uG#	��*X��CqnniOb7/cFpjI{J5#x0w.:��2;����.������)�áG�k{�]�˂ei˵"�V��� �C��UW��A��'�]4��r��c���D0[�ܢ�2�p�/�B �դ�fv�b"�|�>�R��%��jd�}&>�QL!�7��:c��t#~��!�0���m)Д�֟_y�g&Mm@'ݧ$����c�-plm	p�X1}ϻ�)%���Y����1��`�%%���=���.V��$h쩁
 /ө��.�[@�A!;��� C(k��8����W�w}x��h���N/�r�^H���e�-�(o����x��hr�/�0���&�����V�G��n�𷇑Ψx����l7�zքw��K�$�y鿌#ų�>�3�~t����[bc; c�&���04���e��<-V�!J�wAH_*���ZI��`,l�Ԭz&RAn�7�C�SoK/���E���]������/ej3��-���a�&K�"�����U��yۻHR?PWa�~v�?�vg�ڌM i?Օ�AE����t~��hT�C�嬘�������lw�T��<ۥ;�i-�e�M��G�d	�4`=���,����gd#G=_K|2���y�d��
�ӿ�q}������~MX�]�m�d��X��5��g��j��� `-��tF��^�>�<\I�ަY�s�&e}tz���S�',����� �����R�[G�J.E򠢅�Ô���,OkTT��%ha�0�:$�����I����@%X�BG�����4�� ���p��)Sg�m����ݪ�q�+�2��&��kNM[Ҏ1#�U�~���w2��S�I�k�hq5�h&���h[�
� ���|<�ZQI�ǯ?A	�Q��]��c}s�	�L[b�y�a���e,w��D��}��Y���L"�h���f��a j�*��2���kķz
cK°�17qի�vQ��$�K{=��,�D{
����(��R�p}����D�MJu�����?�b���u�%w���>�er@�OC���,ɹ�gKsW_%��1��Z%ư����������F�N��H
Ed��j�'�(���J.K���ȳ��N�e� �tf�4Hvd���ϭ�1����p�)�'+Ҿ�bw�Ȁ\��$�T�ͨ���.��WbW��4�]�l[��:<��C�W�m�O9e�cE�"��}w�K�y�%a+r����!�PB�91%i�a�����e���	X(��?��׆m�������.�\.��!Pw����`�jܛ�,X"G�l��C�q����W������%G��讥1=OӉ�ߝ F�5R2�%,����A�|@��|�6�'�Wϭ������Uu��oW�h�����s��O����0]'��,k�UxF��� u����4FO*8/���$Ϗ����1�Mz���#�C=�i9� ݝ'a��:����^gpK�ˍ��@Z����!�(�����A���Ww{T�44��+J?�2ok\!-A���[E�6�V��/D�o{��m�@��^��s��R�RH �|���|�Va�?���E�@�6�_��Ίȵ��]?:��	z̳@f�C�+�*=)!o��!�\�=_m:��L��!e3Hj�\�~͖o0��q�&Ӣ��O�G��Mo��1Ñ/�i�0e=��ʣ������A.'oX8L��$���	����8:��&�I?Y�ᇷ�x R���A.�7���j�ȂRO\�h��l���UI�۬ż�<� [HJ3���_,�7�1`��>Fu.���
bл��������<?�f�z�N:�!a�i���c8,X
�dħy�]*�az>�(���zw�Eh�(@��6��tR�T�z���?(h��y#���#���HILӻ��_�C�C��U������@bC���Opz.��R�*PY)c��YX�p~����g��;���:�J��4��b�Esr��<� ���ޜ�qA!+#��2���*���E� ���7n��&�%���F�Ή�I��8��#%�0�2���TS��j���Řz�^��W|9 Z���|�ʁ|Yk������Y�grY���A1���|�
s�#ݱ{�(6�J�3��\U�������d����q.�u����d�z!�������֤i�"��>�l�vD=V����֢�RU�WJQ��׺SX�ֱbT����[y1'�Ɯ��i��UDd
�V��ͥZ�?��u��q�~l�{[�0���i4;���`N�l��_���m�ֽ��o�"7�*M'9T$�o)�EZU��S�y����b��ǹ���W2�Xd��l�q%Q�kw�3Da!�,d!�\������
|8�n�x� n���	\w�'h�cU��E�-��9�N ���Z���y8�������o15@����Sq�	 ݭQ�D�N���V�^����-^a���^�x��acuB�H�;��X*�v2�Zih�pl��=���M����Oa�}Ϥ{�0蝠�.UK�_�~O�P�>�ܥ��6�hmp?��QC��6�y�0��ZBٺ�*���0D\��j����%�.�; m���c6s�*> ���2i��&f㠛�v@TD�2u/S�$��1�pϽ��7����#z��2>xW��8�X?����Wx�n���nV�>��i�埙��ؠ2*��}�]��B��2�����>H����t���z����o����L@*�Ī �?$�Ţ/Qm��W�n�A��7sz�gX%�:���6����S��j*�.����zJ ��1�sPG^%Td{-L+���K�Xዦ�v-��A�/��J�aD��8��tD�Eحm�Ok	XU�gI���m��lד�&��;��ݞ�MU�`�.�_�6�K��?_�۳�`Ԛ�L?�_}���J��xͭ�k�.�t�`�圑ݣ@?�V�זPk{�^b?��S�G������{\�A��b�V���¨�ʗT��r�!w2è�LO���[*�*�Y ǽ>d�Czғ;�P�	��X,��^C��7~V�)�4��޳a�m߮+����YXV?C�l#.L��� ���R�z�xq#��<HF���~�aY�8�C
@6�J�&b��Ao�U�hǲ�dX�?{G��I(#�G\&Ei��!����$��HG>F�mP\�̃V��r��>��AQ�P�+J��,�G(Z��ofu<�'�IR���M�Ž�
���i�M:��7������rp�7����ܶ�"s� ^�5ǋ?�,������bp�ǭ��A�����B�Ы�̒eW֡�=��W�)�A�Tk�vs���:��$j��آeL��GH�!��"h�e�Q�jB�]BMA�� ([���]���]��u�2K0��h��X�I��Bz���'��t`�ޤA���1d 
�����S�-� ,��8�J�������4-��X����"T���{�c�{u|��ْ�G*}ѡ�m��pX�����d5_�c�?�W��ښ�X�JP�@���Xa�@&�?��� MO�v
�+,ɎM|Mi���5�)]ˡ�tm� f��3~�9!]�W5�ˏ�9F��$,�  �Q��TΌ��C)��+�Q��,�c+ǋ��ĵֳ��ְ�!\���0
�����U���T��L{p���z0�w�	 >��I>����
�M��Yʋ<�<��fW�{h1�!�CUm��g��j����0���s��4�a��z Z�[}6,{���՟lc�r*�����+�4�K�Z{6Vη�qg� 8��
�� ��G� �Yf؉�|�Ҙ���^UB�o|]wU6�-.��b��L��}yX���<��Q.f����
;�-�DM񳏴8�,������.n���<a�+��������=���'{��$����ڡ�0Dt_r���)�n��ߍ�N�3_�^Los$��VέA�%;� p�*�Nެ�o�m��TE����@Ze��ѧ�E:��D�#�X�G��8�j����r*)�B�$1"��y~m���s����M���䏟W�� Jh6��WA |c���B��y���;G9C$��8b!���x�]5�٣�2-{?����`^�V���BtZ�����o*�↊�t��w��_�hq���f�%�-���'��9��!S˰�%����{Goe����/=�����d<�]|/rzl��N+j����w:-Z�+T���o�oIWy��Jl��f�o��g����J$̆�A��\,uU���R,a��A$������T�1��|Ҭ\LK�;f��0ԓ�kMr���ǫ�������vB�Ct"��Œ곆Ѻt#ݽϫ���!����Y�1��*Z�#V�9��;�\���AkM���҈!M;,�F��| p�T�W�Z��������YKzO��)���VCb��I�0���B8�����IU�HgRr��%	"$H]���ӂc.�h�V�;�k��R��"	a���fMp ]r����~�]��oϵq��^�b��,-{Q�
q|��ytlQ���������S�	�i1ǝS:���5�&em��0�'ሳ���a�x��\[�r��W�-�po(�	栬�6g��".���h��#�qK�ɩ]�����V���`�4����y�#��K1���uGr?�E�v�Fӱ��E�La��k_���ɷ�J�㍸u{^N�j����*�ME���^\�5I�cS��jSQs$�d_�Q�swXdw���vF��=��c��W���;��k�^��[Y:������1���*R�<ɒ��$�>Nl9�ɍ���4���{t�	�+ט��w"Xj��\1.�g�����_)��uCwH�AJ�k�c��I����,�M��7.~{&�ޟ�e^-]k���y���`�E�������8��wk�?�o���ݜi �V�E�T1���h��6��,j_xe!�'O��C6"�ى�5��h�]+w"�����t���[��"�6�
���!_�#�Rֽ��=�Sc ����{M`ꑰE'-�r��t��Ͼ��˦TA�[Ur�[��lm<8`�x/ns��N*���+A,V������ѧ2 �6�,#
mrr��,j�!0B�(6x{��5�Ͽ�`�oHi@�75�"�*+G��d�fqyC+t�8����Q��,���Fz��Ň��5s{����Z�d�t��~_� ����N�X��j'��S(c����H�sp/�Ì��6i1jM`O�G�U���ī���,�h�Vnt;�����+�u�uX��Q0i���_1�h]ت�fd���4$
�IT ��8����M��h#ʂt ��Mѷc�L�`�����W��<������Z��!T��a��l��V5S�8MM��������V$��]'�]ylʀ'�?]��۞+�.�G�-�u�G���S�
/�Z�Һ�c��"�s�`9�uWMթ~*':γ�zG�?�e,QΞ�=|����0�E' ��l�Ɏ&�s+Ҝ��-«�K�EGz,~
[R�}�^��R���^v�O��6�?�T�(���$U�';R	>F���ɍQ��4�X�%�k���m�8Fj����:�/1����.�L˨�`u�߶Q��Y$$���v�-�V�ٶ֋(̪���� ��
�w�����\��ZE¯ji5�0۹/6�p��B�
�f�x�o{{,%<d��Ͽ_ɋ+U�EjFb��"�]�䭌>ڳxǄ����g�{�v6����/F���!{%(C��,�Ha����L��ow���ZՑ�;u�Ր�E�T`7�r�����;����u�������l�e0�WLΨԒJ�b��6�/���rE��KL�&���u���@�Mʑ��`&<9��SVz�1
e�ɶ����	Ԩ���3T9�ij�&�� �]Y�
eB�m���r�v&��[t2&�/�����YP��y�f���c{�<�GH�N��f���ff��`9�|#s��$Z�cW��yr7�H�g��4ABjރW;���^l����V�a�Q`��g�}����[�:��Rў��n�{O��L��T��5)��ݫ��L�ZѶM*��azか���ğ>����ף��r��u{nv8dƕC���
�e��dsA����p��:�9�I�p���Pv$��, ���|��˔�<�$P��4�r+j�2C�k�"a�Ri;f�؊c4��.��cGf�Dޯ.n{͟��vۡ:�D��Cb�M�24`�=f�d�l[	�Ա+�xҥ�0Gs��ʆ�#����*#0=L�}�P�#.��/��Ipń�0����lY��h8��F�E��;�3�%*ڷ��JZ���*���΄��09*�	��wTsـ�nhcA�0:c˧�&�q4J�-��S<�m�'��_T��˶*���Yv5��<vu)�� "�n�����x@�����t�ie��l���`�O�8���,�/�&,�'����&@ġx�N��������(V�%�����M��B�6��G<F�ݍ"V�~׻�J���͟7]�t`9��H�V]�6��j�5���j)���K���6��w%ؓ���q�׈���6�����qr�'j�E7"��gÿe������?��'<�E���)�b�gB%�͗�SՅ<��b����3������d��-󚧪��f΅x��A����Uw�&x��>�/<Ze����?z��{�7�[i�����>��n�����d�w�<*�s`���MË#x��1M�c�H��0S��s���% �+%��z�kb��������Z�g	�W�;+�oέ�=�aR�F�4��p���	�n�PeÁq��	�-�${W��m����ڻ���Ӓ��r� �L;��)�n�]X��מ1�Y����X��X6ٳz0ag:�d�	F���MG��v���Z���t$��p����v-��L�zd�Cs�
J�R�������]p5^�J�Ir��yP��!���j_
؈�K�9�%���Q��0_5���0q���-���F	�t��E����

$-v:L�
�������?O�������
�WBJ�Oؙ5}����)�⑕��&����/l��:���|D9`9r�zQcz_"?(�U~��u��O�ٞ���cIF�����l�I�.�����%��O��s:���%^�r�R)(�p�)L���ZL�.u�{�H���w  R{W�� :�/c`��Q��w�o��F��-)7���ޏ.[��m6w�M�+��خ��i��^��.�y��o�{CzTf�<!'d؍�T��d��~X�rhw���5.��sg��(��1x+�R�O���$����J�a?���a��D||�Ӹh�E��oQ'nո'���i�OEe�r�� ��Ƭ���X4���>g��^������v�5�`���&�M56��G�sq*e	}z���&��v�tdR�	���*`Z�����؞y59�V��Btt�۷{�2��e�q�/�!�q�5b&�'��K�'��m�oݕ��'�����Ƙj�2�Q�v\ >?)�������أη$�KfLm�أ$L�35~��<���*f�z���6�iƋ{������XH'1�*��g��o��L�������0��m�'/��y��8D���YBkt��ʵ��`<4.�@[��l�JʗY���U�w�tx�~��ӌ2�/�q�%X*����&x�������+��8 ̮��?� (X�.��;���;%��'�zg��&��yv�����[�a����04Z9 ��,x��D���४�Ⱥ��-7���krgmDП�B��Im(n���� R�8b�ڽ3�J�|�b{����<m_����Ɉ�*���$�k������Ƿ�`!`,�J��p�'��?�������c�$>���o����j�/?,��}x%iѤup&�c%���~R��8���٫�A�̂�V姚��6j�JWz�y]|���ЌPG+ ���zj�/��N0�Z{�a:q�r��<����#��(耨.'�];��f{x���o_��(�xq�����8��ڞ��xt��~p�3s��*���X_�1f��-��0�X�2}�ʗ�>b�hI�YX"p�Lr��6��1fqP��|h3��" A�� 6���~�f��,�T6`��lt�Dҫ�HJ++��*-�:�]�m���D�|e Z;t_���a!�L���7�
�CѬ�|�d�}p���پ��ڷx��0�vK�r�7���U��kԓ�𽹵�b��UC��B��%��� �J	�c�V�GB7#t�!?6D7�t:EP��gW��f��K0ʶ�j� XǫO/�hF��	+2�kF��=�3GI��7�ؒ�#�Ҟ{�����R=���OΚ�K��]�yyᡊ�Nm������p�{� �:y-!G�M��Z���n۟X9,�0�*��L�I3)2u��^��2�=ut�<l��i/ҡc4;RE�hUģT�V$��s���,=�=e��S~�L
H���5f����k�y>�4�]�P0y�<S���޳+�� ��R���3|[�]rru1���֜x*�9Y�:��h��ì��cE��y}�Z�
h�4q]�5�Z�Ac���<52�zT��G�%>"8>����Qj�h���N�v�y�rt�v;;��G�����P��c��fJ"���|=ыR�u�G��m�w������MS4-�fjt��<\gQ�8TX��:���$&
���Z�Z+R�'L�A����"b/��\y��3@d`U�?4D~�-N<8 pVbA��o�z��:k��p�7��'������%gU�ѵZ�{PY8�؀��Xa6�ͭmsSLU.S>&!6���=db�J�����6
�]����:
���S�l����O"`�-;2��HnM0dv�d�:��>B����a��zy��j_������ic5������ G�vR����C�+�li�A�|��EFVh҅k����jį^c"����G'p���W�I��C?>l�Yb�2W�G�bCF�Ut�E�r6���.5�g���?
�{��;m�)l�J�g�� mp.#�ˤ\�tL�`�.0�I��	��e�NyI�u�_&Ukt����|��������$/Kf��/t��q�{���&�C��c�N�f|@��ܕ�G�>L�ߏ�v;˩Pz��<��_���O/��K� �N�"p�!h*��p�N�7/-w���yX�(����+0�6�|�>n����b�M~�f9��^Q���)6p�͔ɰ��cO�"��b��;��]W�[-�P;�LueV��E8@
��Մ�T�9����U�On��,�� pi�+�*��*%����ⰼ�J?�)��%�]���0UqB x�>n�2�2��}�	�#-�/��������^k�,�<���0�MM]�	���j��{ ��5m+c&��B�գpg`};<��Z֫�XFU
��G� M~4��_>[��"C���2����@��^��ug �����q"��2Ov'WuT�nk�$2�r`^[a�m&�}T�5�Ւ��ɼ�ZQ6lh��d�BW�i}���wYs����M/��\���;���e��>x �Ԇ�FF���\��'�g�|r�\��&T���Q]8����Zc�+&�,#�8����C� 9���a2M��=�&�>�	�\ ��dp��;�p/6W���ps@����s��թ��h��H�J鞙�up^4q�t�+�!����<�}����[�vK,F�&*s24�fK����sq�O�\m�A�0_��dx����zB��-7�n�H�O1]��7,��c�@�T�VI2"�	;M��e����u�i ђ��%�A�vP�1~\l@TT}�Z��5ߙ�g�J%���L�t��S�w���9,��F��΄q8!\#yVW{?��3R����Q�:J��D�"q���F!����,J��"��B >z����S_r�9��(}��ma�9�5�����/�>���+��#^vlK�e������W[�12���]~�M�(�䷮sk���bR�o�0��y�<,�(<��^���yҒ���T+�X�Z鱩�� n��֍z�}�=�љ$Q���F����Uf�is�&4����鵽^ś�}s���Y���F�E��eV��!2��b����
�@��$�b}���g�۾��� ��že6?%0�f=I�GOAe��Oťiu�H1㍦I|�'{77��'����&�̾��0^�Q���<?l�bnyD�⤅0�J}�TUt���s'0�*}oQf/B���}�#BSesؖ1��f�\IN��T5��
�DEW �x�ݙ�J�\����{�WMfu��DK#h��.9����ʭ���n����;�e��ɔT�ul��S[g�ۓ��!�&4j�)����#�ߏ��ML�:nە3�h4$�!�Ynk��Kȝl����	�]��"��_�[+��"�pB��3X?�B?���{�a�RҖ�M�l�z���?��W�T$f�2� (�����:;uN������Ǒؓ6����XAa�!=�zsp�1�L����N
L�<+����w�I�/���/M��Z�hˇ-K�GM˗Q5@X
���AH�#S���܅1����D���b�$��i% �>W�ش�3�6���!�`Y�i2~��`������99��ʠf��+rc���;5t���W��Z��	t�x�N-f�ǎ� �X|Ŏ��KD��l=�W�GE��Q
Sc_�����z����t}�e��G^,J�ZF����t`�L_���:�%�"Kb]�m+ͭ�࠷�>
�W��
5��#��g���c#-̅�#V��6V�t�́�c�*�i�*��E��=�ʱi�Yj�W4�ju^�
L	�Q�Q Fhg#�����;%��tS�I'���$���&��Z�m�����ꥦ�[�9��[f%y|���>-E�W��qJr����bR���`�1�@4�G͊F�?Ǽ��߬�yP��t��m��bDgplFKe� !�����Vh�H�Q���Vf�����7C���^C�yy*�[��|��Aq�G
K�[����1�Kє��7�����d��N�=�?�q�`	��N�9�RT*�D�!�a��R �ӾV���u�Z�ƫ�P�q�L�0��X	�T�xܛ�a�=o��[�i��ǰ�$�Tr����Z�i�*��/<'ТWrͪ$���s���?W�W_���.'��&���@����0����t����0�B��c+R+�0a�A�ȣ����4)9I�i����li&N��*Dr��uUI�,t���4�����To��c�Z-9с�a���Ad]5{����W)�x\�\SlO�ɼ�4~����Yq�?:Fá�`��t���Iҍ4MtZc"H/>�Oɨ&�N��ݎ���r*��u]�R2BoD*��x<Z��B�E�I�19�,�	�N0-/S�T ���L�1��&�Q���f��Z�U�qKn������L2s�Y����u��*3ԔQ�ʐ�EƓ4�5��W�E�˻I]JȈB�Q������i�9}�r�f����}T�Ѱgf��l�ޭ1��*!(�ְ�8�v���
�4��#��I�k�`�p:��ǌ���A�����o�b�� �$�kJ����i�ȁLU#T��޿dP�O��~j���x������SS��:�K�[��*Em$ �".w��ƍl3�O�-��<����	�a�x��gں��xn���5�SN�*=�46�Gn��vO�JHP��@�~g�s�a�4�)&ݑo���kl����O�"�2���m\T����f&#�e�`!�G��]��C�<oy� D�h�!�'N��늶���_ט�,ᘭ6Z!q�/�01�du�.��/�n��>�Ci��$+��܏8��Sz�˘�ڍw��'��`�(��5���I`b�w�҇��pq���XFu���?��S�V�]�����4g�) �i�h���
���`��k,;B��o�f#}���K<"�д�׉lp�ӕ��^!����eNv��r�a#`޶��]{&�!�d������Uh3�)Ӡzf��ٯ�r\�5(cd�	źL�V}V/#	��w�P�&
ny��ӴJ�������LS�,�6�O�8��-���� �x�����dD��J�Ӭ��8������A���_��y��؅�Bq�9��vƬ����R���� ���������n�t}���#�uJ	�<���R�qr���_ݼ��PS3::���h�	�0:��.#��4*N;[������:44蔓�܋}ˬ0l�+|
^^¢������ٮp�1Q���>xJ��v3D>��	M�
e�FLq�z4�.X:��Ŷ(�X|�$c̄���t���y�M˽ Ċ�mQ�eo�a�O�������nw�
�����㶖=��a�J���Os1�����j�Ռ�'ܟN��Y瀻�������2A� ��/���2��?dM�#����tqَH�X�h��6ƢeP�e��X8���i��t%Q(b&Ya s��r���Q��'�Ab�׌�D�J����<�ۏǐ_X��ς���\�l�p�&��n�j����K*���L�z4�U����mz7En9�r2$����
������j���ą@�e��}?	s� �Q��	K��R_�z�h��o����]>]�r���EN��U;6�M7�OƧS(̭p�~�������E9x��AY٪������ �R�1�͸~2\k�$�$RIZr�Lh2�LQ�_JC�5MZ(V"������2З踅�ʵQ:u�?���͕#�,�����U�x��aAWi��^[{X}j�l���c�� W4��vg�|�AES!��%A�]�P��� g受�qь���5�x�����fU6n�|"�����3�	���)����ZLv7���R��X��)��ʢ���$n�X�0�j�x��nI�<��=w_)�;��ڼ~� �P0��9+;�o2�H74��
Ȗ�\�C}�W<?����gW�R.R.�,iaԸ���|q�(!�6մ��8�W���&��R� �gcM���3�ߕ[�,
�$�yU7N�� 儑g���e���E�nM}k'F��$��T�N�8<JɄ�/���g�+���F�0d���y���}ҳH���1���B�$�صOL����^�frVL-�)�R�`�uj�h4�}S��d|�I������˚�ˏ~�dӧ�(���n��tH��b=��	��,���|���
�͚��N����7|�@�#��]��{���HIy=����B`h��r�7y�l�z�/���λԗ|/%�����D�/��E�q<�d2�u�Ԇ2a���$���JH7ņ���-���{��K��)�z)�|kc�:>x-y﮴#�tt�S\$�
���h-�����aƉX�\վ��M|jP���I���_k�Qgz�M��Se=	��2��-~���R��
x��A+���W{>7��=��Y1^������$�-�BV'���	k����e��8|�YF��mMv�A�	;M~%����ٓvMi�!�d>�=�Î����xg�lT�6@ `V�#-��/&� G���O��1��0p	�ά>хWx���ݛ�W ?��>;�F� [�����ҒJvc��LZ6M_Ot������c%9I��K�"��Fh���i�[KV-aMՓ��o����`�ZgM-�jo@������SA����K�%Efa�FF!��=:����DY.?�.�{��R�e����h��������0������Px��NCr�ٲo�)W�s�y
�ٵ�?��r���2ǐی���d4t���;'f��b_��{����QK�D�Ci��c��NZ���T�D�Y��j���-����8���/����
�����`0�P���>������5N��?���޼��I����Z���t@��y޾4��6�|�~}�[1L�u�V<�����A���v\��m�Ӽ�\=�g�c�s��FC�(��. ���M\њ��g�eHSdd+h�f���l���*����{T�=�����'���CI��3��<���&�� ,�^x�(��`���4
��~*:WZ�^�*!�ÞJ&X:��ƥ�0x��=���.4�� G�/t��Ӣ�l^�w`�,6�{� �)�v�=����
����i ���Ki�R]5fQXK^����Z� 2��=���7���#�ׯ���c���#�y.���u���/��"�2�C�L!P���^��=���������|G��«�r���hj۲q�ps8�6JN�V���������Xp��d���8+b���}v\�� ��i%���l�f �{�>4.V^���1S��ӗ��OTwڋ`��ԝ�?����i9�$Ez�9����Ed>K��1k���o��E�w��L"�c��Uɸ�wm�Vծ��5�ƻW�XM0�͑<�Gh@B$jb��*�_�X��{��@�.l��J
F<�_�ACGC����4��)��?g_=�F~\  Yvԍ�N_�2z�Z�hzC��$ȥ��_��$���&���G��?o:�W�&B9�u��;�Wiqf�a�Ҹ�(��g�8������O�ݮ�︝MR^zZ�S��TO��v%`��\Ʊ�dؙ,I{�c(����q��c<[�pѼ�$ &&�X��7���4��[��W��gN�=�)<Y 6��w����u!)_&G�R�of+�e�B|�.���s���xӹ�/2�TQ��=��`�� �<�kR�n�0ޯ�T����:�K:Js,m��(5K`Np����'ڶGW#��������C@���0i��4J��ɕ�鉊����Р������.D�~�^?�nA��^(���d$�|򺑁�0����K3�l�Ͳ~��:�V~��%�ZI�rY4��[=�t�!�� �������	�_��K�c�<Q=��^��|3�i^�O��(���{>K;��3�Da�:H���q;�T)�-�w;�T�Ȯg��!��J�f����i�T��ȳ�er��W��J+4��;�r���*��ǌ~�:��8����Ω��]1��D)��3	m�&$�e���������X�9��O�'Ow2U��e��
,D�/�z�(�K49�����R���o�|��uX�_H��Bm��6/1<g��7EG��'��#Z`��
�2�#��Q��X�k�u!=�|B�c@�������Y��$'_����[�'	�u��^ih�3/���wv)	�9j��y1�Kۜx����T�m��\�)RN�r��=�^_t�[AӴ:hHf�¼�G2H^;�$�Ȍ�Ӱ��Gv1A6m�㡧�Qw B[�d�_�$b-�	���<.��ŀC���@�s�`���V:��k	��Pab@N7_�,j�chk�MU߭-�dw��A�M!����T��n7�����I�l��+X���UH�u;ݧ*���>��w�e��{�Ұ5P����g��M%*`�ȟ������ݱ��fS���c���ʢg�#�Ϥ�k�S�Ӫ���ܤ�|��qd�@�?��W�v@�����vF�b�{�n�	�,�I�n�>L�珮	��y�K(����a1*���2���ҥ�~�2�0F���o~I���Csd�l�(E�����ˡ�3�I_A��NX
ꥶ�8J.��XSuiz�˚b���֎�?zʦ�E�"����wRl8S���3�r��ϫg����(���BE���W�9�Q���g��5��2��l����SPn�o�\Eoย!�ڠ���ڰ;X���/�*�z�����S�3�)������þh��+�)�F�b<���Sl��h�aōF�Ԃ|�s��������3=�'
֑���M�^�KQm�����҃s��+�nߧA�*�^��T������lUQ�:�j��d�&~��,Z7���ݨ��U�������{++��.�h0i�6��>��u��m�M�w���S��B�!�7Nf_2�Q�)���eq6p��q����0N�C���Ϗ$��S�A��8��r�\/�I���h5�-�]�~Uuf�w����@p0)4�r�c�F����pW>}��*S�w���ݺ���%�c���7nC��Rʇ��twO���r��i*1^���C�ߧRC����#��	6�з����A���}h4�����x7������	e�S�i{���~������h(�V^MЎlܹa�C��1���8��^W�_<c�����^+4�"
C�ܹ��74{���#*<aU���]*lݘ��b��1�ළ�WE-se����T�vZ�ǘN�˰}�������ݽX��څ���m�v�A��u�o��1e̴l�,8I
4r�v����"$g�h����W��y��b�`H��@���)�/:˘�;[���S��w�e)��e���;x�K�=eC�i��˥_�������/+w��X�3'&^���i���m�\V�BҢH��;�͇8�m�-��<�˘���j�}1���/��csr{�"s�U+怐���XC��o��P,�i:�|�i�Ƶ!�$��-������`F|B��R��|��ז,sb��R�����9 �Y����ٔ�?	��:�RuFq�!e�sP���N]��_�Bz���}2����u[tB1�j6dy��Ȥ(�Ng�vʾ�LE�h3.3(hE�3�  ������4�h;K�h�(M��qw�:��%�
4��΅���I��9)�I5���>����Jp��\���y����F��sR[��2�RGm�X����@X��=�����E�k� @T�wC��"��৞U���4�8���?-0�7-�Uո�{v�}���Ә[��̓~��w�1���jN��ذd�]���{a_5�2���Og��21���Xp�n�ͣ��7w�[�����:I,����Ͽzt6�޵�<$�
 "���4x��������WWg�\��-Ax��չ�VǪ�Ǚ�kN|���-��nEV�*�P�bS}�3���U�=�B��B��eU���g��=�ZG��/4�QaA�9`93�e��7M�g�$����/n��Ί
#u>#�+�g����g�R�O��T�É�C(_DƩ蜟v�R `Z~��l�����D�����A Z@�p�E:f���[�~Q�-\��#�Ui���)®{���]F=��Լ͔&p����vB����u���W�nu�� C����	�c���aEȾjcF�[��؛�~���j��h�gbt��t��NJ?xC�OSc�K͍8qIТT$`�G���w��ŵ�C��"�p>3ef�>�����d���@������4heĥ�jG�;�oGg�޼�G�������[~�e�R>p��O��e���h�zC��߀���2z�m&}���~�3ۚ\C�nR�1�L絙��	���T�Q�M��ƎF�և�P]�Kc����u+��/��q��h$b�1����_��J����4N-|���܌W4��J|K�i�rf�T�iÄ8^p�=K��{�|�����>s��_*�R��ku��>��u��E��P�<���|���H����zC���]E#��3���e���;.��x�Oe[�������jwC��8��ᨒXOS�{'\z��J���SA��*�U�O,	�/طt~"�GN1�e>5/��b���o�ͻ�G6���[�;$ѐ�9u:����p����B{�4��N���`�%�1t6��,�C�׫Ã:7��T@I�����8/n�r���΢�`9^���n�aU���� ���?%$b3�⯺�1��q��Ӻ_5
WPG�Vկ�_�!��1�������T	��}�;��9��^]�׷��:������D�nK��U`�2��u�[��V-���jR�/]&/j�Vk�Tz�SN���i0����,q��Ipy ��a����5�*�a�Aps86�=�i^�
�ߚm@a'Qh,x	���>l�V��.ہ��2�����GarhU�H/��'F�n����=̚*���F�ۈ	�n��1�
�6�~�r��6W�ʲ!���R�W+�Wv.Y`���<�X��g�2�FB��*&V�6l��òx|9I���7���_CH=���:'��5����m�CX�Wտ�|�k)qv�3��a���Iy\��R��0��Ia�E5����ӵ;c��v�Z�<��k�{��H7L�����jʽ}�M:�!2ܠ_��Jr�3�D���P	�u�Rp�㢊��A@k��ѩ11z(E��:KD�薸�ƻ�.�G֮֡���R��_����!�"�[��r0%O��\l�Ws��	o\�Dܛ� �[�g�����|��-��ZY<UX�kdN�q֕�o�����߿=|��=���������G����r?��H��%s��uf�e�������F���	�*Қ\١��'N�<.J܈!M����(t�Y~�L[�ER���(Ş=�v��%.j��?9*���%N��l���s���̸�BKxZ�"�'˯<_�]��zg�Kv �s��\��n�C��C�G���1i�Y��}��:W��M�F3T�Ţ��UP�"gՌ� `�sv;�i��h�D�=؃��6��&*gb�H�i�)5��Bc�0^ϲ������G����7�S��W�p����}Gxy�N��ஒ�6X/3#VL ��������eu螯�N�����B�G��	�"$L��rȗ��9'��"2��I	���e���a�:�1�ytX[Ҥd�_L~�{.��B�\�Ef2��gF��22?1�5����A����g���(��牠��p�H�����=���V��T9�d���!�;�%�X@=����(MJd�H��<8}��%�� ���	VEs����T3�l���?���F���k��X��w�	=���Z̳�J���M�"')A?���#�R����JI,���y�M�3�b��V�e��}J��3-�`wn4�20�-kP�$%LN��$�=-v|^$ ��g��[�A�5��F�5����B~������6߷��(hXyZ
����Y���K�b� ZG �X���k�:9��?G
Znm�50V�D���<�Zvb�������&�x@��%�z)3x[h`�!W����p6�V�a��.��P1��ڤ�c'7��H�qKᥲ���.�Wq��d�4t�ɏ���_�3h:�: ���A�wԷ^X�k?�E��2�!�P�{_p��F��x/w����6Mef�}��K]���#���b�߃�������T�VȻ"��G�#�A'��g]�r�����	���5Gkhr��q��h\*ҝA�K�O�����w��oTUU��ӤP��k1I��ݐ�&����!�E�c�mW��p��Q�7r�9j���{�Q�}J՟*Qq��1�],�o�Z�)����4��%,�����Pf��j��=���#�L~P��)�k	L�U����<X�!H,1��������yd�b'�d��wC��=�0�o?�~g���+�צ��L�_ɲ��h�}�����׈7�}0�e��A��&�vo�� W�&v�Nɛ����r4[%p�m��Qaq"�K�r�_#:�c�j��E���G�����L
T�M��Pup����cy�
k(�5���t6!~���8}{���>�����*g�=Q[����s�&�ė�/3Q��,,�N�Ϭ�tC��1jJ
*R��'b�M���>YAt\4I6�y���&Ls(G����c�
 a�f�0���V���̉l��ly��tN~N+�w\��6��bAh��v��L�4���T���#�O�k���.(k���Z~պ&׻t�$Z��m(�6GnO)�ٗ\_�_i����x��})?�5m�\��YV��ڐ��pSx:�rU���$ �i�-:U J�2I����b�"�q�4�c8��j���Ԇ��|��� ��(M�(�96�ұ�HQ�.iƨ�E?������Kc/diu�*�ս2̃a�E]�Ti��9��A��h���Z<I���rH^��G��~ �K��A5kEM^��Mq��a��dѶg"s�@���vd�e���7�չaS�Xħw��U(�_g���V+FGW�{�Jq-	4v%8	I��W�l�Ȓ��˸W�_F���G�ov����]��r�,��C�k�'�T��wP�G?x�/Ni	]�O�ʣ/C�B8}�֋�lw}�.��U�V��{��V�Y���=��hR��B7���r�U>sf�X~#8j�����0e�.(�@�\��=YM�m�@�֢|�:f=�Co<VK���9��#&�t�z��S��}���ѳ-U���j5Q}���
Y;E�q� �Q���?�V)��ō����D3w�G��}�@�^X���l�m�<��H��s�CF4gy�]Kŀ| �z-�S���-=
Ǒ�*�.m�_�.æ�#��y�-�'��$'������|ZS�iJK�uqG�7��Y����Eb|Tq4P��IP�@Mpm��a��Hv��Z{�.�����M�N�8eڱ�f-l��o�
��5�h��u+���_�{{�*b��@z�!��RУo]}fA��w�WJR����e��׺�_�T�������)Å���aD����`
���j�0�:S(�Y�Lj
s:�cCu�iwx���{�V�UȆ�	vL��5��d�?|&IZ ��j_F��$��M��i��-�u�fz�g�CfΧ@����z|���6��F@��M)�d��0\ B]�r-�`v�r����#H��Y=�ӓ���D�Z�;[	������d��L��i�7�A�~��a�=�Eˁ2�)��nYG5�F@F:������������w����f��#=���AƜ$x��?_��>���H�\�s+�|Pi�Ts��@�������s��T^`��@g��<S"\�Q��g��o�\r��y�%��T�(!�Vf�����ʇ.�UB+p#��A�/�e��q�֬^OɆ�M�7�Ŷ�})��b�;�$2	���	����̀p���N�8�XU�Z�Q�a-y}T�����/-���#-vڢ/,%z�d���y>!yE�y���a;����d����BB����G���� ;TW��#��^����h�NB�HEI����g~c���;cf.�[�M����yP��.߇�&q3�m�^��}=�~�;8���yABZ�-gc545P����R��{�;��p[���K��:9|@����$3���-�1Q��D`+�5m/.]7�=��EĮ�-Y]%@�^$�9���&.~z��=��9��:n��r[[���p;�C��̣��F�b�V��,�w��tR�ԟ�[(�i:sn�x?k[yU�jkk%4ZdL�}�q�.��c�v3K6Sk�����AȒ6��?�B�r�}���3��m�Q���XfH�~vD�蠟d�*�i��tͩZ��R���N���Y�Q�G��(�W-ꂇ\��"���$��GeHt4�� ���b��s����<�
h�hD�����3".��Tia���Eȉ�X���� �}��f��47s���ݒUtxNh_�<���j7;��w	+���ą{̬�;^v�k"�Bݴ}U܀���Q�5^���
�ڦ��Uq�WF�M��p���|��#����%O����#�g�,�Oi�C�}J�v� (ʊ�����7V�Yv�H�*JRM`8=����u�\�䌪�K�[���M�^�����6H���q�+���^1?{k+DB����c�2b�9�
r�n*tx�����Z%0�6♶���oAݭ�O(ի�RT�L����>b�R�UH��U���
�N�-�^�P]ZD7?����8C���a_Fkܰ��� |ϥHe�J�iK�9ջ,�j�[�[pP� ���a���|�����c
w>�C���&�$ǔ8�Kl����H���7n� ;jMO{�5e����Ͷޅ��ԧzm��q}�Y��]��]gj���f�4�`2#��c@��˶�@�-"�eه� ���ȑ4n�鰧��M�N4xy�+~y�.�6y�^[�S�0^俙���Wi�lꁔ[릉�h����d�����#K*	l�8N�kW�G�Lڷ�E�e�.� ��I����L,����R�Y⇶�A���cd
<�r�����d�	M������ˮ�t�}F��N��βx\D�=��Q��1,�_a:?n״�M��W)gDMZ[�c����	W!m�mJCH&�NP��$�]2�;]�)�h��3E���^x��e�/noW��{�<깶F�K�g�CL>����>�E�Q��&���0�kv3ƃ��gG3��n���t�ߊ��,_h1��ݢ>�,��_6 7�a �����N1��+,fo|���Bo��f�oM�WQ4���}/?'1���#��V^wY��.�Gw������/�0��ߑ�ej�r�H<�N)�'ѢU�#�O 	���ݛy�<�w>�?���y�Lj�����Ϲ��ia/J��Qk˪�a�^M�6[B7�8��אc*��}�E9�M�ֺyXИOUz�S����b��c�����;FP�BoMJ�h�	k�����.n��)x���C��Xs����;��?�<q^�P�c_�)�}����±����d��=�8������iL�kB2���Ө���"�NN�+r.�`B����z�7���i.Uhl��e�Uv"������_e��X�����$s��,�4zD�1���s�gC����a��ONX�d���tƍ�B�.�z[���j���I��$m'��ԣsf��q�{z�8��U�$9D/&L���+�.�t���>��]_�C�!IF9�k�<����{˰�7�}�j-[�{�sH��\4h�����/ѩ���c�3�F�ɠ��¶yG���|��dWQ���'w�$��u�n������͂:�B<i���}��F"�TFr�b�Xn9�.��|��?
�޿�9S��Q��$���j��-�V-.k�@#47�o�팻9�M㋋m4~��W�I�ƫ�����lr����JN��dYkg0K�3�Y��e��@�IZz+����g�!Y�� ��D�#�q���D�,�K�AJp��� ��G��.�f���d.�db����0;�������%��E7+E�� Ƕ����䷩TnѼ"怗���`�Xx�~�c��q�0'���Mۭ�@)��z,�S�XV��LQ~�{�����7���A�ç��
��+�6q�׳���!�)Z���%s��^�Fר��gU[A��4��*�f��nX�MC�3E�����Aj�x�݂�H����;�mŮ�%������4�dx�\���0�.:�.0N���Y~���AH=Y��Z��d�?��(����"h^�"���RDߧZ׻���s�g���]�O�kJ���C��?��'�'lBY��U�4�<���S�7�(��A�DS����y��C`QC:��+ ��KM���&������7�Yثb���9'���_��0������C�һ$<^~������{�Լ*��x�����| �t?d�U�/����'�ƠC:�[v��Ĕ�C�J��q�%E��[����9$z��4�M$6��.D��<~QcvW��O33w�Ml�f����CL�+Ӕ���br�_�Q��$��I�*��,��@@�2z�I�9&
qr�l��+��8�a�:��!c9�U��-��M Km\)p�*uO��G���� �x�s����`W�s�UP�*'�>�y��t�x0�T5ػ|�@�	u\���.U�`�R�7I�1�!:�����]z��@��C,$Q:=b��|z�C�5J!�wJ	Rg�OzjB>{J7���E�\��8rgA?�bGl��hjAO�k5�ED�;^����	�,N�e�vޥ��3�Īrkɕt�|Nl��/hB	
_�x��1���M-�ܲ
��P�X�H4�]�@�I���h��tE��{��l���9_�8"l�TU�OjsO�w-�sد��F�0���m��b�������F���qf�ja�mgC&?@T-���0�K�������eƬ�g��Ɩ��(a�$LE���Ϩ���FV� P/�9��_~K߈]���](�qBb��ⷄ�Y9���+W��l�R/A �UI�l#o�{z,ܗ�g�T�B�� ����#�`�U�s@���\�cz�R�A��f-������B�˷�	�EvK�~�A
��I2k���$	�!����][��%��:ja׬$�HnF��Vq�������K�Ӝ�a�^~H��T$N����n���B^tړ�fU�]�m�@���1�Ⱦ�2�j.9T:�y�.n\4IԢ�F��v��).���[q*�z!|�������Cz��\\i!���YR?��Zג�g�:01�j��$]�f���'V��^�o��xd{	6���k!+g�	h.�	d���c�dx2h�,��:��
��?!�WaV�*qо'8�'�s���Ap�TQ!�i���� Q�����/� ���|�\(��j���y�����Lp�b�KE5$�|��0��ϟ� ��?���֏ne��w�U�����6�������KG>��L���%��F�G���`���`{=�l'o���(�~W�e=S�)SL*Yl�)�M��RYx�E9�`�� �Uwl�ܭ�#z5��Ƅ/����'��Ҏ��ށ�>��ݸ��t�\�܍N]}�0������ف�2?�q��� ���;�S�+a����.��vד����Q�Y6kb�ք�MCB����?��/o�ښ�sډ��-�o�b���7m�􆓟Q��M�?�m���;�>D?z$�U�1��k�*��� Z�tk|��g�>M��ո̾ѭ�J+��2~{ݏ�,��⧻������A�}5̗�,K�]馡1��0|�#w�]XU�V@�u�/�-d�"��ϋ&ѷO�(w����C5������z@���L3��`��`"#D(55�
|B�S�s��2��#���8�Ԍ����%z12�&q�@��PF�ր("7őF��Y��dݤ$��h܅w���0ۡ�. �j�Zp�*M�N�M���{k�21X/jǄz��[�������ǥB��y���"�%�f��������d��*9�/**R����?�0�\�B��|W��h���Z��(t�.��)���]����y��Ԍ�4%۰��tm�IT��v����Y�*�P�����iR��#����!��D[x*�E�a��g�1D��2�r��j&Ɗ���2����3�3y��m���؊Ӧ��P(5�~��K-�`j����Q��>7�pM�Z�)���D���[�����f�'��A�ӗ���Q��4�Ӑ�� ��e]��DB/�ǜCrc5yb���Y�:�'#C*]���-4Q�V`��%�%j�sN=��x���&�w$��h�!ɺ]�����⭇Z��?*M�y���J�O�C#� ���k���C�����7���b��)����/�(�6��s���l�W�e�.�)Ȏ�^Ǔ�"b��Ҥ���;�� \��tl}��~�q�����5�'�^\` ����M]S��cߋD>CPr]+��y0q	�Kd�bE�K���z5��v�@����J���q�"�����P��Ú��8L��)��JmCB'Xq���BJ�9�.]#�SLQ5ЍP��G+�iR3'I0v���Cr������;�󠼫�f����·��Bl~�蕊����<�(c͸�(6��}��I�9��T�"֙�<^5��3""�P`����(�X�ks���LeBE=ջB�O��v�z�u�.J�V�s<��jNz
B/�
�*�l���rZ��+���)�z��P�Qf��%�^�1O =	-���^��d�Ӽ�`,4��*z҃t6�3� ����q����X�F�A$�F]���i�D��������ʗW�&L��$r�=����t�(z��O�ǻ��Ĭ��{ZiΣ��GɄ�8�7M�Jw*��Y�/Z@�j�N�A�OY�E����1N�i�%��C<VL���*��G���x��q���OuQ�; a�p��li�K�Ța�~�U�G�fn�r�� ��2hN�Ʃ�=Z�OR�H��'2�!G��F����=~�y^e����@�q�jb�����<�>���!�_�J��h6*�� �vG)l�zK1��|�i�k./g�	f��Z[c��䣗�����{	��[/ї���.��T���L���	Ռ�@��a�h�r�IF�Q�XR@��G�e���Ac(�����Te��W�q�Ǩd3A^�-��݁gi�ԍK�<�� -L��Nl�Uݣ�l�\CFX�q�e��kv��D`��"T�� :�I�	�B��I�e������@X�U#��`�s�O�)ҮU��豺+�������y9/=�I�"wx��C����)�+{p��s���������� ����l�6�(�r%�l�*[�� ~9̗��^��'�,�T^A�6�[M����}t? ;gZ�6��O����-��"�m�D�	!�QQN5*(�I+��O�<��R�y������E������o���k��N�Ee�n��l�\|K�b�ǼxvP"C�b�]� '&���_W_�ò&Iu%��K	:������d*��+,<"�x~[�Rhމʎ�)�F��y鷝~�u.,��i�2�k���%�ڒ�V;x [�E�$��1X����_�UQH�T^叠�*+��%&��)y)|�vH>w��o��
�eƐPpK�P�(���Q8���YG��w�+���o�6ϩ$٪�zD���Ɓ�4�Iy-g��d�� m�!ؙgtُ����@��%�"�M��mrh�%cr���o���
�����Jz.��V.��{
�G�o��,K��֧�j�}���n��Xnk������%tX��W�=�#�;��j)m�e��,�7S^���t���ϰ)��ofq�x@����@�˗[��X����f�C�dC�zdk���O5z��ÔN��צq�DL�z�g�)��.:���IЭ��ќ����8{I�1�]��H�T�K��n7q�CF �p˛��3��� �)���(�i��r���fS�i�U	��ի7-!
@�CW�Ҍ���0�敆����H�����t�8�Wt��"���| �v7�2�d,�a�U��ŏakW|< �K	z!�E=t<�_��/��{�BoZ�OHB��m��	�;��9��7�ʟI0L)�R@A����#6��S, q�������5�q4��2Oɑ�X��s�7�{��g�G(��z�:�F�����Rjs�w,aV�J��\��-�$�����0�O'���q��U�=��0_�ӆ�Q��sژ��|q�kw�=�q��(��7�um�.�j�����㚁���E.�X�i%ݸўbB� ;�&o{���?����ޯLH�r��+FL��_��|)	7Mc��Z�]�(���{qҞ}S0�A;AnW��gǭ�����-�"J3��~�p"W\����=������}OTLo�r��5K���B16��?���|g�Ѵ�H	�T���D�i��5׼�R��gH��V/���ow~��Wx� }&�K&�d�%�3q	V��i2�w�|y�r���>��[���m�;��x��;����W�?y9���?|ew�E�&���×�����	s�1fݣ��8$�n���Y#Ԃޙ �Uu �k9N���T9P��H�x-:t�{`ױ�z��Mjl�� �7[��`c�m�;~����ͦϦ�{Z'��s:HZ`�Ih��<d筘K��ˇEt>�gf��VU���N�#��g���r��唽 ��]��ry��/�6}p�71:Y�G��+q�9I�NQ����Cn<���K#�����z
0䭿�pfʷ|�n�L/�'�[!9&}I�'�{�97�!T��ՍŤ�B��� 7|���Aƚދ�9)�wV�_r!�R��P������iJ��Ԉ�1�-AJ�����T�%��Q;q&��Z�y�D*^A9���G�GM�]�'@�iq������춉v�~6Ve�WCq%*��:|8�"Ml�)�fħ��o��d���ۧ����ӌ^��sѪ�yb+#�1�u	��Z�2�UӢ�?�O��W���`?��İ��������S�V���w�2wÜO��Z��AǇ2�4�~ʯi��*�c1����,p7Y��@n�u����,���-H,quZC>DJ��� ]��E1iz�aM3�fc@t�U����sl��,��8�5p����r˘0��8S��qW����B�X�����<�!�:��]%tq�dRX�Gxz���	���s�\�"���C�P�Ơ�'�6+m	;/L׊di�,��J�l۷X�M��E�vZ΍Zh;�e��]r�Е�W��g%lI���hW�>��ɕ�_fE���R7�s�*G>ا⏋ܑ��!u*��IG��F߼Tk�������_zZ� 7��ht�I�7t��4*����䁽A�(�̀��P��-a�y�|��\}j\ϊ�L�5}��6��lbէA��"����������ޕ�(�'&�:w���Q#ƕ�#+�,�
��M��C�^m-�8�]�:�}x#�[��������2���3�B\��A��C�:ݏ�F��� �k�R<���|�=ǉ@� �8�#Y6�|og*��l��
�gk�����05�~1]Ҋ�~fJ�f<,��\�l����$��2�܂adYU�;�B��~�ᙵ�ݍ��uU(�j�5�yY6�}�J%dj\O��R�zQܭ2�}���M�"t;[�O��puJN��3<64|��U��Q��?�^Aɵ�
��c�Gw���^br��R�A�Q�]L���� ���,k��4�\��P�_���N1ѽ��gF{9�1�L�,���k�W2
B�P�v��LDnӆ
���{�۷A]��Mߍt��]�t��˜�-ٿ�1D��!�l5�±��'�X�Z�%���-u� 
}�Z�<E�L���C9*<Z�U��R4��4���n�N��m-����}�#5D�<e_�Je���]9����r	�l��\����uo��Vty�����w�b\���e5�?�#�vR��������׸�G;P�ܹ6N�d~�'�T��Kpf��Aø��D�g$����>P�� M����?Y�mΑ�8�Z���sd$	UJ�OV�����"r�*�[��S���w��NW&M���Q�$v6��0g�L7ƽ�=s���GkP%I��Ł1���vM�\;�5�e[�ك��Q�5�ȩuZ$ yZ`G��0y�xeJ�o6�T\������Jޙ���6	���ܒM��W#P ��4�Asd��NԀo�N�#(�
Dڬ�J/d��<D.�D�ۥ�x��+.ny~rbuŻ�Dlu$�@��IEq9�I@R���i��"z����|w�K�Ϗ,�l��VNX[�q�C�uv���0��R��n���ЇҦ���SL��EI�P�b��ӧ�%ZV*W>���R�e���n���ّ�E���4������l��
2��_TA5�E�Hu:`�fӹ���9ee��*"�%RG3���[����l�M0����.t�Ӈ9Ӧ$ۓ���j�|����+����p��Q/aY���v�<?]�*;'�N���x���ӸF�Τ��b֬t1���e��E��}-c���΁Ɣv��5��+yȲ���n�T�FXg�3E3�z�O�%a@�s�u���fe��Cf�
�L��o�E�K ��M3u�u���bo:t���n�춂c>+w75��c����oO��U�"@#�Uz�(��"��d�}c��bl{��I�2A���� }��!�o�@��x:H�\-����nmi*�9+�kU��	����,�@�rm�`�g.NH7G<Ik�w3K�u�.ֱ�J��\"¯�w3 Q�r�ʮ$� \O��I
����r0�%j�����zy���,Y5�n�� �2�M���iQ�u�'vs�p:ӌ� O;�����[����(2M����R�6^4���Zg����)ڑġ�.M�T��I�4�8�A�.�ې6qʷ�I&�R�Y��}W[�m��rh�mt��P�p�y,�^�J]t�2%Ԧ���PM=����4��ѕw�E퇀Yl�' �[��(T�5b�j�짳x�#��E8/���ja�Ooʅ,%&1��6��^�NC����+�o���1729AБ�G�@����8A6�/��o4�H�����1��s
��r�����i�ǁ1�r���f[���T;�����qj�NU���DF����Iy�BX�$�������iO��)
F?��F�+W1����<o�F>�_6�
U�0�{LJsBG>RRb��v#c���q�AF�n䛆R�U��k�:\�JY�|V�[�ӤW��?ۍ�3y͂I�#߂tU�%b��YV�!ye�w<hC���p�l�G"r`�$̻��j�i��<x�@���e���(��c��~;�A��*ر�R�*��|B�NY�ڌ;hW������_r�2����bL�%����8+� Or珔�©��*ήɂA�m�q���1�c�7��
4Z�� ��ϓN݋�*�sv�KJl@K�*Nd�PT���Y퇆w��a|͜ҵ-:}+�=�JWh*����$ü��}�,�z�G�17�l�\A!f| ��,r��3�k����_rh��1��Ԉ�a�PNX`d�T1�� J�0�	��Tr�
zز6�ۄC��S��p��5��W�ѷ܁���z��;��2�o�^[�U)��jV\M<��ǹ{)s����c>��� �\ȉ	&��yDW��'���+��@����Ȥ�����N���"�<�~θsXq�n�CY�Nک7L�B36JAƤO�=�
�̑V!��"����몽��F�{�k�9�'tS����%WSE�A��s��;��D��5.��p��h�{�ؒD�hf\��������v�����e�h^�k@B�/S��2e�f�?��UU�X�ϝ�&R=_�Xo��P��A�y4�]�:�WE]8�2��
I�S�r��%�n������G~�]�/���LA���vzl����8׶�fz}k�}�sQ���	0$]+��H�)��Z���$���S�P��l^H����d��.ULt���cEv#�)k-�>��� ц�1f�dU,ѣ������Cv{T��f���g��,^�rS|d��r�̔�e˾j�0z���9&�� �r/ό���Z4�a�F�$IR:�R�T��//��կS�B�l.������sj�K}�쯀�b��nH
�w[٢��f^���\��� ߽mH��QI ���H�u�Hr�Z��ې�~���1��X��W�&5��r���C��	�[�#���-c��wӋ���D��U�p͛��%234��x�Q�mQ����o�gP�
���Y��Y���Y	~(�y�i�=x#���6}Ԓ%�����n1�����͞f�h)Η�Ex�`uO�n"1��vh2���8��c������J׎�R ��C�����3��>�F{C1S��)��90W�"���IG")��U���'U<�ɲ5�շFo�T7 �B6v%I���]d�E��o3�����I.uɟ!SlY�>w) J,�l���+7x�L��z�W�'�{0��-� �Z,֯�J)%;baGN�N�I��;���fGA	���ѭ5:(!^��T�}VŦZ�O��䧠RA  ���<R�_����vh��p"���&��@���ZX�P�Ⱥ{>�=���n�ZZ<B^�<�y�7�M���^�n	ƨ ��P R*!RO#f�>�[�ʹX���N��J�Z�����s���u5XR��mcV�u#�}w�H�f�q����W�8f[!o	�È��:T��8w�+��rO��v��h��6�4;���>'y�^��ERLҟ�a�m<��Td��9]��?3���n.���(����K֌j:��(��ġJ;;�{�Ep����n�'Y��h;�[QDč��O	O\c=�����<��ں{��@�V��Ԅ΀�����LS�B�[�!�2�=�y�w��
+'�[�nw<=�%!�EZ�}w��4 O�qN�~��+DD�'{�N����*Fjb����R�+�08��a2�D��aa<�`�~,��m�I[�h���FH��b>u��瓆	UEv�Eq�[̒�O9��z*�I|�aq�� p�T��E	�y3ƿ��J[�q�6(:G�&�w���C(��OR����]}"ϒ޵�A):�D��j�ɷ��&�je9H��f�-e���v]Aow�1����~�M�)JG�zy�vK\V���=nځDhd�)�Jq�g��I�1����cR�
�.�������äk~�<r3�.y4u(��Y�՛"�TR�(>��9N8n;�&��b����
I��pN��H�'8N��L(��5�C�e���Jd���xљ
�"<�W߅;��7I��xߠ�Dmc@rr�����W����*�2��"�y�*��p����R"3�D>�٭�D7m;��=a����l�!��!�qjXB�f���ᇼfq�ȝ6�[GDT�P�ӏIR�7x�<�QJI���̙��$�7!k�$��2y��z2�֗��zuR�������(,E��B�$D�`��L��iJ��l�B�sAm�~�n �6��f`�&*���"����Y��97����M��Hڧ�QF�z���߫+���?��_)dk���ޝ)�MnT�,��eX��3��<m�k�B����`IV�o�~�DzB<���L>��7�K�ؙ�ц%|��V�I��Z�r�Ob��	X�v������{Hǽ���dB� r�qCS��-ŏl����e�C�#$��y�"����u���Mmo7����� G$��}�<�#��t��-ۅ����ms,o�a��9���,��r:+�Q��xC��o3?�+T7�R[L>���z\�%R���̑d��ql�I���YXC�V���n��%k���H����R�U��s��"��ʬŴ�qG�L�@�>�q�"Z���ߜ�}8%�9/n��`�V][�݈�J{$�!?o�7�)߼v��N�%�9�ZS��CYG}���ue�M�L���a;�(c�B��0m��G��	�m☡P����ˁ<�����k.��k��%�w�!�~���!!@&�X�0Nv����B�˅.!�����|$%���r�H��(M�r�������|����K.��a� �����z��6.�~��,�C�=\Sۿ[�J�MR��Ԯ��OL�O:^f\��6,�>"�1� ��AH�
��c8���ឺ���n�
���Mت1 ^��rv�&3f�^�jfŪ�[�Wy����d�Z��*�>����=�����M	�IGd�0$|n��۪V;�رA7�}0Bte��hħ����܄!��N�؅X�� �k�9�9v'�.#Y��z����쮢}�OrM��H���L\��߉@��3PR���pfr��ߖBu�fY�"��@쨘�y�N��� ��x�A�ki�z�uk�<���[*CfWל�4g�����)��z�	uL}PE����he��ĳޝ���|�=<%�rT��>�I>�JE��#R�ձK��u��7�0�=�*�C�к� :�-���(���<�"k/W|v���>MTݘV�!�+0��� [՛�v$���6�z�>�\-Q�g��C���?0|XP�`�y�=m5��Wt).���i��;$�WqSfY�T �>~�d>��R_��i��I������a���M�X��kH9a�`ܿ�#=�I�ڈ�~"x�1-,-t_�8��1�T�n
���ҫ��:yc��i�W�ݓ�צ�Ll7��>C��A�'���:XH�M.�7��{r��P֐�����,$S^�>bXK5�qӅ�Gc�Xj�%6�8?���J�jt{�A�?OT�X��h�W��Qav[dC85
A��3Ɵ ܫ}AjSqp''�(`��4C>x������NO!�	ZiN�Ĕ9��c"k��<��'K��i��qq'�����ʹ�Ƽ(r"�!ƍ8�D��aި^�|�K��a�]���V�9��3�*�����݈6�r� ���?���o��O&�Q�l�ĐV���\	��{o��Yeti$�bt4� JE���5����l�o~g�{4�b���6�����h�}4AAi?���'���;�t�-ނ��o�&���mdB_wZNNЌv8����������i�k���H9�]����V��}f��FJ�O�Oޣ�I�"dA����Ȑu^s�K�GXZX@���:(	,���>1O��Mkb���Y��Y�����*[N����P�8�O�z]�n[�Ba�?�+*w�*?��'��L��Ӵ�Ɂ��FE�V�3�@�:�v�z��pF�)�zsNg,a�UF~E���v8��g��u�?|o�c��P�(�
��ԣgvx��9�X(������%�!7�����2�Xb��E!{�:$����� �/��cO����d�(��C�Δ�N�\����)��w��	_>础��f�)Yl~ŭڿ�(������(2.��̫J�>�M����x����C�~(���}b�{���ɂ+pB
�8$��� ;'�q�GoY���G�F*�'�<�$"���)��ةHM�F��C1�,����}߾��t��Y�"�g�A�	0l�w���|	x_�?�w(Igw:"V�Zj��0��0P|T�LU2��^,�Ҹ�/�%ɑ�b��������rA)�-�&dd?�Cp�]�P����eGYT+���zE�|S4�+����&?��6���6��FPJ7-�әԬ��}�ao�wfc�{Eл�3����˧FC�BG����w�Q���6�Ed]k�ao��ۛ�dǟ�#M*���n2��Is�*�U����Rö˩T5m1������S&ͥ�yn���	J)5��L2L��o~��@��m4d�쒹Z���U���	`�k����7�Oʓ����׵��X9�a�pJ��@޾y��§�<Ԧ������h��T ���B�$���R���=�&|�91i[^�ə�T�o	����h-��F�{�쥛�՘Z�GW�"X�^˕���F������{;���bR�;c����Y�c�&�w4_K�T�����jC7�z+Zf�#�i
��r�m�>bv�ms�¬k�Hñ�P��!�����p-D������A�7��J��y��� s�3����r��Nå�����|M`�˚��ݏZ�C1N����@3^}T�|�vVH I
"?8���r}z�fԽǫ�ٍ��x������9�.��(���)�t��$��ƽ>��͓��s�4��hV��>}�jb�T7ּ0����R�17.��Ϧ��n*����.� �E������� ���Z��i-��*�U�����p�E��N8���NQJw����KV�������Ҫ�e���� �OQ'�˨����.�%%=Uv98!�T}�.;��Vl��Ijz��TџW	MY����:�کD�wŊ
mh�z� � c����LE㪬b���l�X�m�έτ��r�F@��I�_���l�:� 
�w=����$�
1�ȴ�'���;Ƌ��9�� BM�w��������.xZ�2}
��(����R��oS(�F�����������?�UP��s�x��i�T�r�m��9�b9J�%q��,��&�l�DV��5���$K�^laQk~R �V@�A�E��P�3p�Xv�Ӭ#6�<Hb�c��yu��$��)�dU	��=JH�k$۬ʚ�ă�B��29���Q��[]�z �M���c,�G��H����3��rT|�5��<�6��GRȵ�3�#��P�zEn5���M^�DłK�����^�&�ɗ���$_!ޭ"�qv&�켄�;�z�6(� �e�
��+�I7����ML�!׵d vf,[wT���]8�Y�G+Տ���m�_�-�/G�	̀9�f��IjDV�����=�8Zѱ��=�o�R�����m�-V���X���fTTn���T���Y(l�b�C��$;�.Jl}�b1��IZ�G\=�D����S�D���W%�~���tqb����[�S	=��u�<8�x��(m�����٦��:��i�&Ѿ"�U�1�	�qn;�]�.�^ˮ(6�Kb�|{Z�����!z�)��.�=��$ @σ� n��㥞;�����=�$Bp��'x/���؋1��i�k���m���7;���8������ӎK+��N�o�TM����TxbP��^�PGw�G�5��N���1���O�払��uS��J��Q�X��I5<�Ӄ��,�0��,P�C��h�ߛh>�*ÚLO}���2����^x�{�F%ʶi��q��a�ݤ��?��6�,W��}HS�D�f��z��/E('��BL>�9!X.� Jv����(̲�w#?�PZ�ľA�'6�:�G-'Ͱ��d-퉠��{_�0o�tˬI�E[gm���j��;�	(D��!#���4��|eT�@l���
/�&�["��xb�o��(��Cע�2d@�?����S�M�=��窐u��E�6�f�.ֶ�ȫ�)�n�$�^O�P�ϣ�~�{�C����!��5��*� ��7�qs�0\T�����wK��a�U�G�P�p����x�rXq}�dm)��XE�E�c�<��0g<r@O�i�ژl������t9�F@M�}8z�H�Hzp�1�t�ʋ$��_���/1��,�I!�e�6����������w��{��"� ��F��sp1�9t��e�ԯ.�t��Jo��&�X����o�d��4����C?�����+q����Y�����`����VUpƩD&]��<�x� (��i���$�[#�e�ߐ�2Ts��q�gȾL@0$�ZU7�����G�?*J;�����5|2�9�q@`|Mq��+�b��L����u~��p�#�l��D���_��[��I��Wt�Q���w���h%2P�3#TCt����3*Vc�:�z��{+�a�q{k���q�5����J���ߕ~��D��(��!�S�
��k���$i!�(�^�Y&L��ҭ	a��s6  htZ�N�66�n�kq�����Iv�%DA��V=�A����
�&,�BX�k~�m��E5ά��5�@�ߺ"�9�߯�
�-6�A2&-uȲsb��Q�CC�
u7e"#�L(���|��i-:7-�7^�]?�Th;Z ^�[��e\��j�kۮ���*@f6y`��&�L�	����WV�(*��T���3_-Ӎ ���'��COP�fn����F\ڭ��M����9X��(���Y���B�9T�ŃDbU2���8EMb_��HM(f4|����x�N����$˔O�BI��aîJ
�F�����7���l�d8�X�Շ�v�����!�e���vZ���+���&��YƢ����1�<�]o� �Ȗ{ǋ�b�6BQrY�H!K�b[~�+���+V��H����:��Z�]}��������h��!�!�fr��wt?���^�$U��Ml8<V��!�z�J����ʗ���nN�2��(H��K^��2��3��b�gM~w��=m��t�KG���~� ���y��I�'�+�4xӾ�B�h��]F��^7EWܑ�Ka�y�W}Gy ���	n�Nۖ�H#�O�|�o|5/�� �N��[��l��%�v)i,M���Q���	���!�er2m����S�_�4�d�f�@�������?��-�5���~`W���cfÈ�����P��K�ܞ�2\����d!�<��kR�Nc+!b��Y�1g���y����0�6$�4g>����K|��SC���>���K��)3k�Ǚ[��P����LէV��pt8�Lo��1/,Α������8�΍�.mi#/�0<�|`����]D��Hk�[�p6= W��NG�2
�\�%�P�h��}�C�{C�3��R�{�͟a4�m�Llʻ��ܜ����RG���|%���f�Ψ��T[�u����nj�+ÿv]�v���򎤂~y)5E��~���ߒ q�_�XXs_o�C���˺ ;\�
���٪���d�3��H�����7���Z�k(�U(D��/�g";��-�~Up���4�J�N_w���R�FA���2�}w��vD𐦂�ѽ��A�J�C���"���
�aGV���^���SA;s����t����%Z#i8i?=�
��/;��kE�ש����+�Ԣ̷h���������L���	w{�a@���N�F¤��=z���˃ϕ��YI浤B&�� [¸����++k1)�D�H�%�4H�}�\���բ���.2�߁��f���a+y��[4]��Q��o����"\�Mr�|�y7�� E�i�f���6���̐�E���h�p3:۞��&��׃���F����W취���<��	�)�EԔ�)�&�Z��8)��in2I��=�y8���6�^%H��]}�pT�����I��}2��z��VXܽ���4�5��G�F Bd����6��'�t.7�}�e���'���Y�D�iO��EI�������Y���������W{dW�)E!7�d^��f�="d��̝��
m��=Caz�<Q{эD +�βb"�#Acv[DH�Ay������#���P>��k9�xX�/���f��T���:q{\w��Y��9�ˮ�X��:��I3 %Ϥu{�&�z�deD7�1�8Kߖ����>��!}��dG W����r����B$+{����x�߱2�����x���(q�����Q ��\[{�A~mԷ�Ci�yfƗ?�;�6���T!Wl8ݽAO%� uC��4��k�"�UXq��`�<M��+���+�ۋˍ�U��V��f!�:��ۈ9u��T�|IPA�@��RCk �n4MƉzx�Y�T��yw����+Z��[(����d㒾	V,��T�U���:x��	��#2o�y^��;���4��b��0t�mA��DHX��g�L�Wyl�ˁ A��c����]��aإg�n������q����	&�Bsf����Cɴ45�Joc �V:�A_�F��*�Z�<l@��bB��Y������^�p7%��6�"���_I1�$4�44s���~� �9��I<�J�!�4���GI��oopvxNꞗ�ͨ�iAQ9iD�
�{ {��\�$`���Q88|��%j��.��'	Zo3�5ʋU|�8��e(�M�M"І�Z0�p�C�1�$� ���j��I|f�oVv�����vXH���Vs���|B&M�:���sT��o�h�JJf�<�A��)z/���̸��&��|zf�;M*��/��v,�Iצ	���N���ا���Ve�GcdT��lK���Gq��_��h�uX�m]f�@��?��q��Y��u�G.l�%E��+VAwڏ��q��凈q��I9 U;x����S�BY9rzQ��W�����n��:J�z�i���G8 :*�]|�o4@����˾�M��ZlY�Q�f���
������(~�=<��w�~=2ˊM�8ԕy�K�'����������R�y���S4��������w��8��͸�m�E�Z��X�h�B-g&W��5�i���t0E��H[ux�W�a��:@�s*�� ��	O�����ʶe���f�M�2�/dxHY+�a0/�C��4U�3�iwPQ�(�;	]TCэ���]&�O��!x~Bfw�< ���Gj#AN%���C��$�e
(u�wl�'��L_�w�n߀cc�z����N� �u�7�C�/`2=����HN����+]��m
2i2�§��_�Ѭ�Cإ�7ă�>����'�>G���/ y��-:j~.3��C���9���\�w�C��<��/��
�8Pg����#���~�������1�䦎+#�M߷6�8^�O�(���	>�m��w������st��uu�5È|u|�0p��W"Hخt2����������0 �M6�kkU�A�����f���C,���ƅ?��Zks8�VF7^��\���ں��]�bn/?��R�xN&���w���s��sy�;׸�UvM�Z�|:o�{i}��'a���U2��^s�ۊ�&X'$E7ԅ�Ϗ����A&��P�
��"�ً���������m�$i��*�ن�����J����ilX����	�ݞ��_c5�LI�TF�R��'y�(�3lܑ�'Y�<� �b��d#�xr6�(��t~_"4�Xo�DO����_I����Ֆ��&w;���1!s�I�e:o�bm�W�4/�7������L��J�*����m���,��_����7������?����*����h�>jr�,�c�I��\>���DhI����M���ұ"{o:n��ph��%���,qTG�T"ha'�OG�x�����&S@�J�U�{���ؔ�Իg Sت��x�F/�uޤ*�F��d�<�Y�Rj�
�㢫���w�S����`���D@o���f�vLE�ɏCba��9�g���r���%��<�ͣ�/���96tl�^l�h���w+��%YA�;�����Y�M�7��M�;�x	�ø�00�C�[�,��뛏�WDuN��&�aU�I�����2z;7�{2�sJ��޹T*w�\�?�yZ�d~�C��1h��.L���C�L|���xܹ���8��?e�h�6*��Ы�S���;Sn".�Qs��wX
R+b7�Ժݷr�`X���9Yᐧ��j���m����0�';��K*+��F�d7z�B]�\,,�j��ǤE�[`�%�KqI{A�SfP���%.9m�e	���m�)u���S�o�[���e�gb���D��uT�G�t
h�ca	�mi����6��!�T4�16�2H�]<�8z�w��������Gs2�LH�f��l7� Z[iP8<[��q����`��BiȈzq�!惟Be�R���f��`3GZ�mk�|�;6WqVrYQ���A�8�O�жd�q,3�#�y����{��[�#I�(j#��4awpn`�n�ո�l�x��38���ع�w?U��5���l�;`��f��6�4=�n�SO2���qk��S֬�c(��:��$�����!��K{Nt�<����|��e�+�Q�?�
�l��m�3�J;N���R �hֱbkSWG߽��H���Ō|k|<P�|��EYo$n�Ou2���zs�B ~�X4�>*h����=��K��iK�ҧ�_��B|�$�[��gRR߰s�j�3���-��sN����B����Y4;$
�'���`A(��y2�A!��x>������F%��#�"�B��%��u��v�e�)��/��>�SĻ����$�n
˔��u�.S����]L�@��m�$H������bw�A�v }Wd �$��"�ᅠN^ͱ����$�L�����my�ށ��]�������߽3AёA��f����ԯ<gp��dWX�r�ѫ,��o�+����KeTVBOu��c1�7�{�>m6��Vvҷ���B/S+p��Y	T��/+�"�lC>�N��5"��
���2�-�B��.Ğ��Q�cp��#K�s)��%���|�0��:��q2���u�����U���prK��}�!�o����v�[s����S��u%�m^�����)NXd}c��wG�\�>�zS��?&% 5!+�����Y���	�{�=�Ul-�\h�9��N��&�����%�4ef�r����igwo]e�k�%9��6+{���{'�!���o*:��z���G��Dw�<��$����9q�:lOiӿ\�bW��#Yo8r悔>K���"ZX ~��a���@}��bjd`qfFF-�rdxL��NXV&�z��g^K\?����8�L�:����d3;O`�1�I�څ�zH�/�芾"�T�~��¥��!�n�N	�hA��S�����D�)z;�Y�ly�ƌ�@�j]�1ǝ��?���0�ͼ�jkb{��fL3r�#g^!�>1��X�x�iB�LhØ�*p8��]c����|�ؒ�gq���I��ʹ��{V��š�9�_�ӄӣ�L�+蜷����kjF���d�k���r��!"+�/��0&���"d�Ya��E���Q��O`T�#����獋�݆�)��lF��錖����ti�Y*��� �%e�5ǣ��C�����\��Y�e��i�S�}�y���	!�RiO͙,L�s_E��q�����Z,�*G
�Td�-�t���$���ţ���j�=u1*#�,��<i��_��S�wk|TsL��S��fV�.�c�107�O6k��>�/�D�\���&FΫ�X���� ���Qd��nM��tU�?ńz`eE�իSM�\�"d� v3KU�?k+m=`��{����Ů$|jP�+�y��ţ�=��u��1�ط�����B��sB�R�l�υ���}�P,fgvw����;��Ofa��=H�LZ;[-�=�QG�4�G%8�y'��wM׹nʛ.�&�q:'��G|��GNc�!*�2���Y�+��T�b��v��6<�K���c��
-ނD#V]�a O���*�h�s8�k2(��"ɛ]��{��%�p7M�W>��&Ar�W.@�K�l���vrS��C<fU�l{ �c���E�E�,���sk�kۻ�j�I��ؕ��L�a`Qn��fg=�Tĥ�,_�*�@��-��D��KD��b���x9bsw�f�$R��K'�r��	�)�\@��X��J�p��=`�:��|v�KI2���z���W��k��Ni�,�/��Q~0"�tU�M1��1Y��`��s��\�t�@�~E��cR��)W�>��J0�H"���	�]V�C�௷L���XX�O�&r�JC3�`e�Sv��a�מ/gӄ��J��J�i���y�x����)(2_�rYL�����E�C��B�Ư�!�C��G/j@G�t0�R���v���%8���Z��˪ �§)�cy��M�d��(�hB�.D���� ��&�&��25�&��(����Y�����B��T*�V���(����d���VP\��{���ل�i0�e���I?�X�Ь��"LI�6�+��ޘ�8��u�b�@�q��f��m^<������}p��h���(>�Qg�E+��� ��}X����X@��+�J��Ħ��tݚyN�$BO�u�Z�d���O�X�2���\ �����������*� Z^����E��2����Qr\���~�*Doh�\pOc��r���Mi�*�cg>�K�J��л�2y���˱�BqF��W�`�;DO��D/(�1c)�B��F��F��2� ���2�ʄ�XW�H�.V��z%�&�w'���`P�K�c�ic�r����^�f�"��X:,>@��ٯԡ|)�n�]bH�C�~c
�3���5$S0�K��
���,��Lq���~�
V�ji�#B�u�2��7ȫ/"� ����v��F\T�s��4�MP�c������l���S���)��3~$`od���e'.y;���-�F\��B��D1���L��N��w�?��
��u�ZWTb���H���&$��u��_m��'2�a��5`Z�ٷKv�j'妦C1̎��W�7�#���ɜ��]�j�wO��r�e-�Y��`�1$m�ږ<�^>�4�~�����"��U��d%ߖ��6�,�/�۶EQT��fa�,���w�A�7mI�)o��oB�k��ڴF�� Ty_�v[��W��&J�z��`��/2b2+Yh�G#���;c�Da�P�u�A&��g�V��b?�bJ���/��w�i�ɡ�)I�!M�k��u�k:�=g��������⧊j�f].�W�oTn�7������:>�;o`����������,ݸ}�n�mʦ��!��~��6]>\���9`��yȈ�4��lѭL�� �����&�/�0G���ېrl"�p����x�ܿ�1*/SG5�G���h
o�V ���J{(˼���dJ;kNǌ�h�֣iu\��k�����@�vՐ��N�H��J��碩�KP�V;x�*�p�]�ءHX>��AQ|�΄�`�:���(�������j�$�?���:��k�U�	��e���ʾ��,�rbq�<E�ie�R������_��	�8
Ӳ�D��{;������;s
��c���-Må��\eoS�A��v���+�\��{�����ۦ�.*�𜩣��Kb��W	�k*d7j*wC��p�Q��r��Pp(��4�VsI�!���d~1��F��H�"�ʄ}�\TO�B���n2�ꇀ� �G���S��ْ,�S�� ���V!�'ių�g���A��Lj
��kd4R:?����4w����/�M�g�g�/X��P���&L�����mwr޷R�DP�Fq����8�O5��p�6�K;���\g(F��E� ˭�
�Ϧ����H��I����vc�r7���� �4G��e�¡���`�m����'z_=�΍ؠ��B�(|�f�|�gB�� eϼ��s��V�{�r*bq�ZB��w�i�qy៷ՇX�=e�������B/�@@o
X���!�Fo�f9�G��_v'�m]:Y�����P;�+���>ҍ(������N�fFt�0�_�����O�	}'7 ���U�o Ϝ��馩ϝ�열���˔uZ�C,r��v7���
<�LP�5g���~�+m+�X��`dB��'�����kQ{����bpQ����9
U��[_��U�-�u���Ј���y~��-�1��B�8u}oW�zJ�~��r��QGM�,�Z�d,UE9T ��+	ȲF�*��AS�ߤ��\fX�mV[cFB�J�]v����C���R��V}�`� '�*��@�WS�����O�� �i)ʚ�pV�A���wy˜vd���T�U��^�W>�{݇��.2#�TN���4i���Qrʕe�8W`��᠆����Y���k��bm>�J!��#��v��b��a��GT2�̰����#Z8yӀSb	���5�g��dz=�@	C���|������{��R�����*�#!����*{LO���|����F�ve���
�3'ԙ!�k���Ŕ͇�R�N���*���kst���&�X�e+
r�iCq1^�)jb᯦OxY�}��OD5{!��62�BJ}�֘<�@�ǥ�m�j��ƛ�·�xS�>=Yd�q���u�s��,�Ӈ˖�;>��o����#�]�P��,I�R��PcJptX �֑Y�Zj�_�*���ɶp/���_� ���s�<�z�s�i��=��:>$�m��k���;��2�ڳ��P=r�u֜T�����<eߎ�8)�=�ނeӀ@����f�݈����^7XqJu�|%�-j����"�q�B���K40G���x�@�b�z+D&�8�9r'�J�n��Z���������.��)Ƀ����P�#��QYLO�;gHxg^�n� �R�f��@��I##2	����!ʫ�
v|�dAp��������l��vß��F'bO��8�A?�l�^����kR���HZx���(A��@��b:�>)�ەV~ҵݞ�Co�a�Z!W�S���3���O�͂�eD��GGh5P�G�F*�� P��&�[w��@�����%����K�Cb^������!�x)y�u[O2����J�J9^~,Wt�&x��zK��9�m���z���p�k��{�[
q�e�n:�/@;�P���etɶ#`D� ���51���*H>'�'J̇�}�+�U���l�#J)ǫ��Z�r��Q-t0O���l�O�- �Z"��=I:��&[^)Z0�:,�������7�_#8P�߁OCd��=:��@��Q�2�>�S�(I?iut"$�
�-6���j��	kޝ�*XG4dd��?�6�Fc����9�a�X?�<+�,R��i �K��7Ѣ��>B�E߽0�7ק��pq4D�z�XmKI\
JȲ<J���,�c{9)"�Z�=$*¯�(I_�L��`�"��	�8L��>��q������˝E�a��֖xm橋"i�C��P�klb���G�3�I��O%K�&�M��U)�e�D����ŷ+j��+,d�ܘ��K�{_lRۛ�>���z�����'&���d��3Ҳ;a#� �{�
��4�H�Z/-����\�]y���&I>6��7�8o*��+��;�ܿ�`�%G!⫏�=�Պ�U�?�:x;9,Hd:lB�?Wd��HM�*������P�VZ��*b�i��U�V<�o���r�JC~���{��]��a���o�4>��D�"8��<���#�8���D7&C��ov��|-�������#1��ҡ4��"�aU�5�jC'ȼ�_�w���b��K�����h��Dw�6u�~w�bW�q������qt���oϟ��`��<�03Sy��!��7,��վ��$����9�N#�ꃹնu�`xD�<��Dnt���G���p_��9�u� ը%\4�[f�9���z��:O��E]���K��l�V���R���/��d���b����)�!^��-$Er/ i:������P�C�G�#���E�������V�S����8���*���X*=��8u�Y�nv�N�y�,�q����s��pu��2�)��Y���ա!,[�M�"$��	wޫ�m�|���:��������?����
w"č-��m
�k��It�viec��Ύ�gP��^���~F�g�;L�=&�Ss8uO
��y�&��_���۴^Cq�Y�6�J�
;6ᯠi5��ѻ�ލ��M��SAz3�������okn8\$P��(����W��H���Tw��S�����f�4�+SLq��7N<�|6��~���F}����n�F�4��ΰJ��q�j�o���.�=�;�ݏ(?��<������)��v���F�j`6��C:'g|G�0V�n�*-��2���_���P�b�H?�~�bG����f��f�Q���%��¦'�[�T�W���ԥ]��u���ј(������/�E�B�\桕�?�E�s���{o���ͥN]N����8�}(-�H��r�6¸��= ie	��#�R�0��>�V�	�լ����)�fz�"�W&T������I�g������Ž�:�rb��TX�`���r���ɪ��Pi����f�Њ����O	]:?�r�G�	�y7���!���T���9A�C�?>�&j��F���;!�bM��"p՘b�c��MLS�3�������,���Ab���oZx1����R�S���6�����)�<����20E0����T�6���H��< ��Eܠ���V�ԆiT�P%�?�~��>�"�+����`�K�������\4�x�x}��g-��B�f�H�)�b�e� >.:"}̮A.�v*$�����n�g]����~�턴"] g�oS��
�r�cE����y��d!�ڮ	\��6�;+�͊x�Xa2�r�U�LND����� ��{�O�p|vՅ���L �Lp!�R[m7c�Ґ�T�\�h��dv+.�^c���7O���(�|X�j�ߊ�dꎠq�S˕��(�<�{�čmP�������H׻�HO�L��~T}�O"X�?�p�{���ng��aC��hD $]�	?���_�I�D��al��N"��p����ur����W���q�e�p~�ӓI��F@�|}v��h=�!�x~�y�E��'�'5	�6��R�o�{��*>2֓J���Yx/���*�hB�}�����ߖ�o����j��E����sf�e?a`�b�t	j�\e�4&%�B�� �\Y�s؉�J6�h��"�>���[��b�_y����-�c�sO�|�Ռ����
���o��gp��'t�%�װ���j�W%�U�M͆pK�
w_���I��x
vf�b?� d�^F��e|.����@rS?� �F�3 ��i�x3�d4��v䋇��G*F�i7��z�~ ���Z�r�pҎ�H�w�(P�h^	�^x��xX�2E�_�������V�=Ɉ0g{�z��D"��(���g��J"�ln{D`5g�w�d\��0�D���Z�� D[+x/�{4IqP�E�H�0%P7i2Ì� 	G�S����	�D'u")=���]t����=�z ��(���A���eG����W�Gz�r�);�+�o�g��X'U;�zjÑ�1o�,�Yq�f�\`�]b�6[�5vc��y����\�-ϋ�T���h;�j�*��������3�<�%wξy�7iy|����g����}"gڶ����`��9�NT+/�3��~�	n�b�2���ǌG+\0	�\��zz`����oﵫ��*��#���7�o>� A��;X#O"gL��y��l�E̵Vm��a�J��騘9�]���K��9f�xR��䢢I���+�r����p�铝m�N�'�A'M�߂�L	�7qA/~����T�{�q?�@������=I{�7�:�B������ᯍ�0*V�~f��S��/�"�>ꕘ	^��)��I����#8���*��޿!pa�b�|a����9��&ZgЇ��n�(�t���,-�]�wa���'y�W+�M�Ħwy�����}#Д�3��F j��2즀��P�@M{�6�K�<y����E�(�VO�#��.z�'�* �omD��nÔ�|o�B�DW�	�L�}��(�}H"��1C�-H�����h�ߩ4�O#,i��h�#BV��t���PTw��\�^1ݨK��2T�jf��̭:���Gv�%�E�@�����X+Sw���(��G�xm��~�;u�=�)[�`�e������q�Y<H�=�x�M�����	��܍���ϋ����O��֋�q�C�W���`��	TCIH)�b\x@�$�V���1�a*H���(CI��)D!XWB<�l_�a&��e�A�����!�����k ��:��D^�?�0{�S'߫�	��қoA{ތ�,'W�r�s�K�9���T�����v��AH`eI��y+0=H�[#�@е��?Ɍ�:��j52����/Ԁ������;Ǵ�Ҹ�C�l��.��a)y"�d �Ӛ�E����D����Z}&et_{~�`�A$�el����8��"���k�:�-È`t�Q���r���I��M,��l�J�H�GxE�G��B�x�S� OBw�|h�y�;�`�O�ī��=׵���F���.2���ϦBL��:/���#��T'�±Gn�e1Yu%6}�������j�>�i���xe0��3�ʅߍ�w$z�k���/4x���]s�r�s����,���"+���p�/ٰ�'}F s]�a����=pkQ L��M��֛���tdxk�|m��9�D<��=֔*r<&��5M?7;!�k&�Ɔ�����k,�9�ŧ5=�K]zi�t�Et��],��-��m�%���X|���k�8���Cp<�{��/�}]t0�*�ry�S�xJKM��ӌY�sB���`�kV��19���,�Po��7h�jd�W�w@���c֟�w���y�=�:c�8lhc�+{aOI(�x.�¦���І{f��{��t����3��Rq�����Xw۷�Ԩ�9���d^ku�G"�5�=%�9K�-�u��gY��]�_�g]��>��GWg'�w3�������@+hf�x��*Ċ�T���	y�?7!�5��V��/��\����rP�cO��>�9>��x[L�Jl1�tӻ,3aK�D}N�[�;k=*�;q�'){[��3넨��9��hQ�kT�_<��i�K�2��^C�1 ��ؠ��~ ����7��i��|�yH�v��$��nN��,��7���/����v��'RWʅ���&7CM����
�`�k�-0ʹH���u��^כ��]�y���[nh��$�t��E��@�������|�FK�pU�<� ��5�)�Ii��&�34'�J_!�sxgu�� �`Ɣ�����/�����O��O��H;�P��&N����`���t����-[���(�zSq�bV��sO���Bm�T�H�iR��w�]��2�\��e�bb�盕ϡ4-��:qS���>8���p����7ֱw�~�ӒA^�'uv<�m�X����isE(���4�#��ht'��g=b��n7{"_�|����Z�2����7C�͍h��[�ꛧcO�GO�j!)sp�i�ȵ�ɶ�✜���N)�Ǝf�Q�MV�����%���3�>����%j��^�d�������@����;E�h��o�����]{9�2�r���O`���y�s	��%e�P�tG@5�l�@�Ko�1䤇���jPaGql����t��qm}�\�t�K�7���vt͚5��ܓ���MI��\�=OE�>�SN�3hS.\�'��6v�M�S1J;/13Q��d�7�S�n��������ȷP���>��[	j��Ll	����ڹ䆲������Fc)����M�Ǩ��:��+��Yg�!u	�a�[~�m�'���1Fza�& �q���v�s�y�'�	�H�3�4�u�C��[�ἱ��O]��w~�|�S��	�IMI�~Fg��0�U'�ɷ�M"�n����z�<N�3��6�����d��gGE��u8���O3�6�W3B>����a^J0��x4�Ir�Y�v�Y,�z����v��&�#�%R����&�TgV�K�x ���_d�S�(����M!x���:�BW���3�����TW3��s�2�3���5�~��;Ҝ��A!���%0�������i���7>Ij��`�J��l��j$~	|q79�.������`�P���H�Kg��C�Gq&E���
��K��ʸ��(��N5qK��r�G���Ak�dgǸ�E�Z��Q2n'��;I��ͧb�.O%%�0�ē��T�l6^���=����_�uZ��jkw�86�� ��^�J�Rc8�M��]��l��,���ì$��M27n�T7��d!�!�o��ᯄ�_*$=��q%r�S���Џ���l��?j��μ]�6��A���w�
@�P]��ޣ��4�׻�	7�B����$/����Hn�B�G�O�x���dOfı�^� �"MT�̨�(t�6ב6�M�E���.��=s7�&���v�����H�忙1��������xO��:m�-����"�`S(��~&S�gq��d����b�p�d�X�E�
��V}]F�L��9�?J鰈��DrHy2�f�#Z�y5���R'Mkp`��_]x?���ÍT�w��
ԇx�Z6{�3�!?)=6*�@�+�p8|�Ȥ�Ͽ�pg���'N�q0��<h�W��Y���j�M.2Գ1�cʹ-.�LW�9�3��n���14}��#��%�M�N���g��%��G�xɛ�nS��+��͕��zl�3��~�2jf��:��̱�S��"��QX����/j(����ӪN��f�0����4۟J�|ۻ�f��:�z�x{� �h�SR8 ����Ja��}�Q�eA,��E9�����"G��E��f*d�>��@�D�x���0Z9E��o��9ߠ����2�M�K񆻌�j���ȀS4s�?h.��|�@���:�t�h���úO�Fp�ˡTG2l�ݸH`hU�~���2�e��:{�h1H�p��|�~)��T�"D�("E2��7wk�C3
�
AѸ~��C����7R����YF ���o変��ej���9��/I�J�4�7y����j����B�����1	!���;��O���Kdes)���m)��ǐD}L ��᢮xa���u;��a��b�d�p�q`Yk,�T�c�ؔ��T�
����i��Ɖ����������ս�b��~�UG��-�tX�����%źxI��� e��ׂ;��O"��v��NI�B�#���D��#�B�lFr���R�Ϥ���Q�&�4Mb��2���o(�����ֹ_4�5u���hwA�E��nDF��\�f@|���dHЮ��OE�gS�@�O#S܂����%������7�Wp���ٕ-If$W���6�lݙ.���(�.�}T'¥�k:bo\~�t�p|����!Nq؆���EoH1��H���������\H�}�e٧�F��`���G3����B����ќH��.�!��)1�mj�[i_��>YԵ���o��Ý(nG*x~�`&&M�D����"31�`F�L+�.�R5q;����:���=rT$BG�7N��괃=Z��H��ZaY�o?��x�C;���Ů����7�"a�����*zI��V�y����-�7 opL[{����R����.��+9%�k�ԟݯ�jY<,�@����⻌V4�7�T]���5����*�b!��
���)�ԇP!�	H�ASo�R���$��T!��ԕ��y9��
V���&=��i8�y�ɞ%\]���7���^d4)�/*A�q�=����)Ƥ����A�B9��%u}rS���U7��2j5���9�vﾖ���Ro(�)�����޺?���A��D�����n�یR��T�j%�@PT�mB
HwҥF(H��_2��f9z����Q:���t+����?��[Kû+$}���8���x"�"��~-�-�ElI��6a��)�,��w�u��:ʑ�5���]�Al��4�<�ȇ�ϑ��l��h�m����cu��P�HsC��Ҹ
a'
�!�j�^����wnԅ�Ӌ��%�񪕻����"A��9 E�xҟ�����`Y��f�E��)�&�f��7ٙ(�0n0)\O ��8�)�@ƒ\zA`�&�u��=��Od�ؿ��oֺk�42$����ܓ4��������A�
�i����9,`�p�n}\�2���*�ѲךW�Vw�~<���Ͻ���Sw`���@�?gJ5{tez��Z�
YG=��~��ۚAp����}bQ����՞�k_8&x8}��ߴ��.k��FJ��ږk�O�[>W���09.�ݨma:��zoV�+Ds��h���D�7��	��B��q���yߚ��(1�P��Q��kPu��[:�"��pSn���ԡ������B�#~��CG�?A��	x��w� �H��o�a1�3�˶��g�[�q����y}6_!)��u[9ޜ�@洌��u5#�A����`�2g�ֵ߾$����S��~�禃�����-�a�K3+=c�rLT�c�w�y �!Jz㧾��D���R�@p(Ip��~��\��X�؅���ø%���|���cI��@Ü+�a0p�W2��m�{���'�?��m�nA��e��q���@2�H�Q����e ��0bA��JI����ꂱB��Bi�ӉA��u9u6�~�����,!V2ވ�P����Z-Psv�,�~ƭOq�$�і�I�U���Q*���T�~����� 0I�	��\|̾`l��'O��3�9�tGb*$x28�Ր��
�7-8�?�aڬ�1�f_���	��I�@���"Ø2��}�r��?Q�C4<�}�RX����eOtҝ�� zd0>/�q��lU�� �*g-�l�M������}�ܗ{���w����E.Ы�4����(3`�{��q�B��DU��fan��O�#�[۝���(���wdR�	-�5�Y�o��������yf���h��ת��2�Dh���Zг������\{�\V/�r�5����,�.=4l�xN,QD�f� ��3X��	B�i
�T��?
��f���|�����d�� ��t�́a��.+a �,V	QH	��;E�:�ߟ<c�<r��<}�ş��
:�Ѿ4�
&�l���?��م��B�v��Wd��ùU�n��Ћ��ώwu����2��&�������dВ�fQ/9��&j����H4 �җ(�������Tf�T��&���k��D��~����dא�y��#��ɦ�v�aq�'�nd��bq��!�S�Q��cm|�W��}u�(HV��߂��cg{��u�i3q�\��w�$��~"��v��2��W�	���G'��4�خ�		�C��H\s��`����w� �N-��(�9mn�5o3zE^�A��*z{&�t@��	Sd��ز���4�i�`Q/2�H�De�x#��j$�׎c�U�?֗�Y�d�x;!DW�������A(]C��e7�1j8a�$�#�v�I�h�I*L��큜�J�ƽ�ʩ��i�ɬ���ӂ�=U���J;X�v}3����E�N��ӃQL(/�糨�)W�kl�U��.�5��>�I�#���z��89���O��j�ވ:S��l�O��W���	�D���������B����`'֥�@Ĥ�Lc�TT���%}O�+�Vϣ{�/�y��Ay������ٙd��ؒ��('�}�o���������%��S���~�VC�&_�y(�i���,g��.6d1���Y:ۦwPK9���Uz)�䢖����S'�_�N��"����6iѬ$��蕙�hx����w���{
4(K�J���Y�)ބh�;�[��X������0ߣ�?v�%�2��|QS��x�����5����l�Ȁ�8L�@�ڮa} �]v�cRѹ��%�#kQ�����}Y�4���T�#�1'���ϱ=D�t������u.p�E}��~�K���U���q?:�u$�h��׶�1 OܲU|/�.(����E����on�3���#�5��m�kF7�-XPFS�^2�?
���a#�2����B��О�A����-�\�k]C_��4
�i�8*ԧ4z�*I3��Ȼ5��� ���/����a�x��y�$�1��ʷKp7�F,�:�Bes)4_��.y���0���΋����ꋣ�{�\-h��MI9��U#_C�����W���d���9c���n��mLړ��!ʃ�Č�|��l��!�7�BK	y��oV�r�נo-^H;oX��!Z�4�
���ʹ�����k��Z� �-�.�R���Һ./&3�ѕ۷r��f���Ƥ>�%B����0e��FD-�ݕ��{,p�2�y9E�,p���5�Ý�u
K�D+��8H\:�0y��sJeu�D�g��/K��R���٘f�Z����*�z7��o�(F�aCT@�Q�`�o�v�����ua�m૝�ڧ��MC�x�����y��Uc���s��
�T-�^
:�a�P�G�\�5{XM�+8������3yD"��i���(�1���h;��5פ�9^"��p#�0����xd6���,�����lk�#���	��ظ%��"�㋐߱�e�p�ݻ�/��Xh(
ȂZ��gp���#-���k=�c���|�y�k�E����&PF�Oz����������N�v��/j�0Q�!�"y�w;PT���A���|��r�����؄j��t�ECo�x��	��ʞ��@5�Zsy�Q��#�]Pc��#�3���6v����f<��aR�b�4�<�#O�F��el��d�Aig�����w���bt]s(��g}�T5�s:�'-��
Nއ�R�I#CM��X[��Ƿ��y?�{,B�51F�#�iƅx��8�z��4��c�M�Q�bH���V&��m�y5���y�,S9��1��:E�5��A�s�9�=uC��	]��ͭF�'��m;���b`�����P%�Y4���:����z��ơ�̟�h�W^���s/=S�sQ���2T�#ަ�ޑv�t^SS�Z\��RU���v��z��>�{;\��w��+�k���ts��6;� W��B&�٫���^�ic[���C0�e9����E��xZ�������1�6��<���
D��|��~x���T{�4yěU�C�\�o)�z�6��)��sNXݺ�I���9�Mۚ�q⯀f�$�lmZ�)ST �G�e��T��ɼ���=��^�%h�i�ͨ��Ž�����һQn�v'�F���:ϴ+����9P1�޾�2Ġ^�V�@��Gf�yX��?��7<ӹ���A}���k��b�{v#l�,d�wh@3�
�b�{lu��Q�aȆ��8�p=/h �Ɛ�c�x-��C)���w�_VtsI��B��Wo�Ӑ��v3f�A�
���/.d��슍���88���,����ޕ|�F�ٝ{sR/�妁��/��þ�Kٕ�=�$1��_�%��vQn����pj "k�������8&���64�ܕ��ݞo'�EJ4	?�; �!��*9���/q�5��f�o|mc�Z�C��z,6gYf<c_��{�k��wt�x�����퍍�vC�o����\�v9�xp�g�j���EW��h"a�RC�E����T�(�Kh�S.���<�G���v E�	"�>�Ӥ�>��6SIQ@b��KN�u޻���n�-��
.�msa}(6��CG�Sg�x�4�!p�l>}��;�cPt���98���F�h#�����YS��2m�pY4P�Tx�c\���)][4U}X9:���/�t��߂(��iJn�Ϊɯ_�gA ��EU+Ȥm��������)bh�C��,�H�نBcp	�M��X[$�L��_�����z�; }_{�tй��g.�Ikf�_s�H㌀O<�(���X���]>EU楞H���gOYAD^���p;��~����S�K���Xg�7>��w�n0n,0���4���kp�GLOtb�b
Q�b�
�]�5�-`:7U��Ʉ�=m�d-�?�֖J��Ή�3��:�i��+P�<�u�cf�SMW�n�I$��� �"�Ϯ�2ܔBZD9nT��[	�2�R1�_��~�)���=�4�6q����3O*\��a[%����$��h׏O�ؓ��&�t8�狂��{5EN������O��1H���%�L��%8]H��[������T��K�U�DM>�O��eQ�!#:��+[�
v���(�V���Q?�DO�?p�"�!�	V<,�jކ���`շ�gz��=d6nZ��'<;�{���i�����>�R[yo/E,�}N��Z/��͙+���#�B���U�YjTC�ē�O��µo'`#�U5Bf8��b_ .��&����.����Q�R2J��B򥙫��0�-�8�?؏@�R��t�O0�]���_e�%��؏��pZ��%S@p<Z�}�h��)n�i(~R�r�_���o`	�H�l@��u^���8aȷ�=y��}���Ҫ�\&��n?,QF�6�F�J�\m�=�x�!��>��uz�z���;���$��r>ծt�;�>��dm�mjy~�L�Y�V<0�]�0��x�7�3�mD'B؞+sb4� ���%N��)�D$X��x��}(?�m��A{qT�}�I
8V[3��ߠR�jh�D2aV#���ũ��Jg��
���㈝D��b�:�Ts<��Y�R�@�(%BF����Q�j�c+�������b�������,�����)�!��aHs�����Ձ+�#�ծ�#�j�T�	_��z]��)�;A�?���&�E�V�l��rMt�����ʇ^�1��7ϻ'aA9�l�S��X�j ��K*~>'n�d�rn7|�?v#���;9?fQW���2�rŁ+aw��_�e�Ӛ��.�&`L�;;6�̨g�n�'��YE�wꍹX;=���@ȟ>���hr ��?Wrx�=~��%T����B�܌�H��N�&���g�S���S�]D�wl�C�&�\����>هN��(��a)xQABf�Y[����cyO�1�w�]9Z� ��}O*��
��i��&��z��f���}	�B�ИM�SI͠����J-;����)RY�"�L��BB|��~S�^g�Jx�$��:�7�'���ON���L�٩���깟����xњX�E��A��4�F���m;����$�6T����&ғv�JUD��6�A�Q	�M<<��p�D�%GPE.T	Ǔ"}.9)c�6���UIJ^������T~2jF��B)�Bԭ/|�IWG�$Q���)������yj&���/
�6lԚnt+k*�K$xѺ�f�V<h�1��}4	?���ĝ����ٻo�V���O6�8#U��/J�����c�8��+�M�U��ڜ貴�g�)���ҹQ���b� p0b�/���-^y��;��ւvck��_��8�8�z���fZ�?�v裘�g���}��T�%����p�:���BSgE}���O̰,��!��x'9T��6�vD�oRH�[(d��F����t]a�4Bd��M96k갓�����N �u�f[N�҄������������9y����{n�ҭ�N@��=o9�Ae 
-�?vD���
|O�[����N���@�۸&�*{X�e=~H�x�Q����j��Z����k���!�G#�	'*�>���t�;���Zt �扨vJ\�1-�ޚR��/Q���;3pI���HJ[�@�EI�����3d�M���p&-�rh<���D��F���nvW˄���g��(��)6+	�l�pB-�'k���g�a���%�J9�Q\������푂��{�y}���c1���I���˳�T�m����Q���s����իM��}���E��O�gjƞ���[ݥ�_ϭ�M��V�4��niZن��  �(2BӪ�6<� ���'mSNI+����W1c�� �;I����������Q��o �K���;�'
\�=UQ|[PlG0��Cp㖆�%F�2�5�>6�O;5_�U�� ��-����t�Ù1����_�
�ε��bA/��4^�C���TM�,����@�&�V\e���v��QM��i����j������E���a�It*��]o���v�>xU���E�x���W@[Xɟ� ������.+�1�;�
B'IG�^�sQ5���+�gK� S����Mm��-k���`�0��n��[,�E�V�h�/�5V�mi� ,��9���k�5R��ɂBxC�P>�Q�a :8�ύS)�|��j�.��,�Iv`���7.�K+>s�����*�@��Զ���@�q�CN�t��:n7@.ƿ�͞�t�I9д���Cs�<y�X^�"6�N��{����s�|CW���AV���#>�2����P�	�f%�QI�}ҙ�7QӁE�>: >��b��
���p��ǈ�����e���5�RM����h�~�� @b�o�J�*�yb_c�++>o��%Io舸;Tr�IQ�+K�,�F��Ѱ�~��ġL���oT�`�E
3��ô��q�YtQ�����~�6f��YWqYK�	�7Z'�홳�n	����'�ot��Y���``�wX���y �Y.��xi�Ұ/��h���ZDv�_�:��	�4�޵�����V���R

��j�E.�&ݖ� }��"<�N�h�AO|]�ʋH�Xk	�*��'���q�_�TOf�C�O�ٷ�(��R[Q�b�@��F)�K\	�����*�B��� ٽ��@�e఍^�Q��a�0hf"�9\i)Uv�V�S�@���h�8�ޱ��l�^q�wY>OO~��(/$wqp-��mX1(��sڿ"��s��¯v�]0=r�N�3�a�|S�y��>2&k��b��Zn3�uKE�̤[�)\9��+ɳ?:R����K�j��r��e�8�>01�����Rr���S�K:蛘p��Еtun��r��I��!�^b��4�dq��v�0�;�ܢiFƯ-�q�EO������_`ڕ���Ytk˓]���o%
Dm����Q1'^]�(�#g|8_��'�*��UG~њ@�qЎB����w��iq���	�1d5Po�:�)�V�t���뫃���Yeĵ乫Sf��U�R���|�9݊�A֋��U���`'������<��Y;T�?��A!Iom��3A�����ꧥOʔ�p�A!�?9l�+�U�-��o'4f�#RD@��v��XC�ژ�%��A���'t�pi�[�8�y��b��!TI�$�Տ��g��r9���=��c��؎�֜3�c�ĻB�ި��cB�"�߾11�N�'�ĻC����wY�'v1��*6&u����$y��A�K��y�b�l�伝)��a�JV�m�uھ .+��C�J�ܽ���t��CG�H���ǻx�ꞚI�e6|(�	U��
B�S���fHE��rq�	�ȗ����J�P��9��Z�����K2M��p0Pí/*��'*���mr��@�sUHk�sj�����p�0���Řf���;�:�=,j�Qh�A���"E ��4��c�hv�Q�z�&�V Nɦ���{A�e�!���"���*:C�1;*�M��*tش	is
C��Lom�A��9C%$J�b!cE���m#�d8	_�%0�F�i/8�\��l@�'��\�����K[F�퐯��O��K�`ݷ+��s��(>g#�9�x�S��6�ۍ��/
*߳�xθ���l�7XZ��q������%E�Ƌ~��2���R��O��f
~<@$ ��ފH�C��D'_)�Ɍ-�{��+�j��᎒pZ��+c�E&��Y5j��c���1����	��G�߱�$�@8�X��b�i���6�����P>�֙�>�P���}s��i)��~����CL�8J�h%�e���yX)�f)r:N ^m��o ���e���S/I��ͱ��%��x,���8��Yaī��m{�h+>�d���e� B�裾
r&�Y5�Q���{>n�Ji���.�Q�VA��*q�N��J��bC��ADo?S��������.3\��|���q��^�:U�xu��h���s��M큱��ęA��I���^�3�8i�1��|��e��wP�a`㋎&�����{��.�	�՘@$Z@{��#X�U���u�u�Z
�Hn��@�wqkC@�ڎ����C��X���;��?r��%�yq�ω�Z啹�j�z��D����"�����D��߹��F@m����oNGTF&�R�W��J�-�� t9߷|j���f�6�"������H��eT�xM�0��ƕj�r��t�R&�����Q6������-���x�;���<hD���.�ik�7�a~�L%�Ȫ�K��`t�B� �1+�z�Si�w?�m���p6�,����D�H7HQӓ�fOk�[
 r�C��iو��z�U��~JU�y7�m�c>�R޽پ�˯�e�����'A<�~��VVa���6���q�٫�zxZ�~b;?ޠ�&{����T*s�&so��p��>fpV��}��x�;iP�bH���i,�G����Q�*=�F:�}g�Jh	G*m���I�M2|_�gQ��j�����+-{��F^�0��B��������	�L<hQ�8V��z�Rk�#Y�Tw�K���pY��N~�"�����i�34&ѽ��v���@�i?���l���K|0]�;X9}S�_b��;����\>��a���<G"w
�-������]ۜ���(]��0?Ԡ��z4K�a��nz`���еz;U�	���I�ֈ����呑���e`�X��C��邽ZÁ���"1�\wr���Z�������M<R;�xV�﫭�d7>E5D�|(i��=���ߴ�� '�c���$̕$���S�� ȑ/1��u1"�'�ħ�k�a�	zXA�;��� ��eȯ�R�Q�}�Κ��A��^!tC�\�c+W� ��}R��!��ׁ$�F��"�}D")�7 y�{� ������c.�K~_�G  �[?D�1Va�ߑ��:��kp�ў�憜0Qi����]�� �CK�m�+$�򻑖f���.ƌ
mx�|t�P��^+�k.� �dn>}9sg�ӈG#7�]�fT���v�Ud�aL@�u�r/5���5R�og�����\�y�6]�Ut���4���9RNxY���Z{�������b�\�쮙���]��:&E#��35n���۽|�a�4��k��/g{{d:�iP�׌e�t�R��tgg������8V��h�&�w�a�q>p{H�Ւ��hG�H{��h(��H>�g��"�}���9(�~��UD��/!��k�c&=�`����&�O�d.�<��6�&²~�H�"ay�dX�Rvpd�N��{����f7u� (�oYULMw7dg��kGz-�~�X��잞���%�'Y��;�1E���2���=,�CM���5�>�S�P�^*��~6'�8��0&�1u���ַ ��H��;�^����T)�uP�O��r���f���|���&6Q��i����*F����$�~.u��Ƕ|k�q_�_@�N��2;5*�����[�|�.=��ˉ+t;��qar�>�u��(W�-��iO�3�C�n=�+`��,�8��2�l���@3���S��i���'%]y���i-�\&�%��$�А ����?��X�����������F�Դ��@h�oP
-P�z
�Y��n����{>	����|/�P�2f��\��j��*2��ۻ�!�>Te^�&�N��}ʄٲ���L����4,��
\�n<�cUS����^ͳ{��o$��!ۢRLPRBm�/��χ]eDk �v뿕;�/��o.:Q�3%N�����I�?ed%�������kyj A�ԓuBC��V��5ʹ1R.���Z,#�3�歋MH_%���^���*u {A��b&��%HJ�?�J�3 g�.��p,_)�@�ͺ�8Rp�(?��;S�I@10	��8��k5f�H�n!���k�ك"4�~�~u�aMx�FSQ%a��8y��lgiܟ�жy�G�N������ĒN��Π�����<��]BI�g*��Y2�C6쳐��=���g�2"�׏I��N�8���{���6��������{�<�Y��}������EXPځ̢F��%t�''z���;>]�t�A�a�_�%�%�9��v
�����W$DǾ�JR��G�J���(u(�a�qEۼ��(;�[�7���x�'F��^��9i凾���޵�'o�Y��ӡ[�j	d�P
_�(?�յ����n���*v���Su�FK5�#ĳ2�i��~�Sp�3����	�I�����͖��3����i�t'p6��Rf/�|y�<��D��n���=%J�/�������3P��B���k�n,���4��������c�pr�
M�L�p�ل���f�g�������"�ps��>�����R���J�;��#����KY]�Cb���s�Ƭ�z��3�)-�d^��\b�9|J8�����,���I��p�&�����Yħg��k��Pe��.⚰ޓy� �e��BT�28����=�я�Iz5R�,�-qW�����Yo<�61�b�a�r�ud��-��7 ��{�.��"!��B�/FtO��"[�h���x�b�g�46�p�� ���%dy=V���vi��yC��a��������($��g��{��K�-�B:tj�T��RNI6+�N)clf�Hť���&���5��94��]�0�	��Q���JO/Xqk��G�$?x��!/|��.�H�=Nv���Y�VN9�+���I���Bs[
�:>bb�ML-,��bۗ- ��ʨ�F�v	!ke�[����-Y�����'�8Y�~'��S7&�z.ڊ�_{�Ϝ6KoUt���,pH�d���l 쪁7���.��� ��ecb ������)������Hª��˴���<���� ݴ9�6-XW��X!c�ZH_����eO�.����$N{`�<�����zc/�p���|�?h�O��a@Ꭳ&��"�?K-*j�8�i�_�Q[45�A�Ѡ>&WX�#=C�T�UL�q�����U���[Ή����0& Yp�?a����%W����69��k�<�k���E���sbI !���E(uB5�K�"U&�%Z�<DE�z��͜��D��8T<�l�d�h��ڤ�;"�-3n�赊<�+ݴ���J�u�R�<˭�3Qo9��G]�������!��I�������:�DK��=+!��m�˞��"�4Fɝ��^Di(��eo�9���q��D�ҩ!BV�1D�%G	�*�j�����>쯄�t29�)�����-b��7,>���k��9�L*��b�D]7��	��<q�P�n�&���^��*߯x,�S�N}�	���434Jg��c��.(uZ@��kt�WOr�4�>�;c�?z�P�tWъ<���ȴ+�4�&{DX<���� �N^؉�k���H�Y�kj�[����U��k�`��Av�;E�0�$��:��ϛ�@,}V�qGh�eG�m����IZ�1u](�zo���7බ�����f��u&��������H�1BJ�`�7N��抠�7=�ܿ>����Iقx���L�]lwOr�H +6�n�E�<� �3�WE�#��Ȧz蟈e�\:��#O��Vx�݇x�>�uX�U�&��'����s9.B7�Z�`�\L#)���f�g��-�LY���kt$k��څ�O�s�����y w� �9"��-��2�0���y��:n�\�Ҥ`�#�+8j��%yf4�~�t� I)��F$�CO�^0�dd4,��o��h�0��_���8R��I�r	G��1}�s�k3+%�l�V���X�-��G)��E�^��j�q�b{�e$?H��F���tV��ϭX�/�6�E`���z�:�ԗ���D���'k��h]�0^K�$�Y5�2J%
r����bd[&��
�&x|�p���{�7e:?`x8u��-y0�sQ�{q�w`�˟B�"�5�ǳ�~R���N��~�4^-I��PN�aԡ(��1��$�"���K5��(��3����:�FwK��#R�{��m^���Mȗ$�
6=9k�J0�oc� ��^8�7�Z)ɽ����KW@��`��^��4\*�-����P	}���ۜ5��p�p�B�9�	�W
�^��A�Jƿ���R�e���`l]�h��{[ɔ^H�p�.�$0$%���!Qn��9���P0��<�k30��R9c/�� ��&�;��=��[�8q����\���q��Y��$Z�a�!�~X]#�uh��P�G��R�EyI��x~~��ϳ�����cM]�'zZ�U~3����h9�;��ԝ95�^�0�6|���V�n!�U�<%�ԙ����4�Fj�_���0����\���̳oL�+Z��^�ˮ�^Maƹ��S��Z��P��)2+��3���̗�6!t�5��i�?�	�%���ß%�o�ȞqD��E�v���m�ƆQ$�{�����ZB��<ۮ01ܖk���NCU�H��5���?�@��?��$V����us�L���7/2�G� [Ѯ� �m7��͡O�������~�%9f�`cۿv2�뎸����a+`�2�W����.^���)G�;z�3�T�w���Ϛ�enDgO�U,�33��_�����/
��'�a��"�4��'1:�_��Fʨ�!��ҟ8+��G����s[�mi>l��v��2������2T��Q��{u����q���Z�w^��3�&�%Gw��Nl�,����:6/���B���3��k�PD2�^��L��0&oZ�,�а_�N�T����0aРc��X��K9��/{��1\ܡ��eЭ���{3)~���D��v�5�~QD��<%D�c�Hd���Ck�](:W�׳�Q�2�y?nW�H��C���Mݝ���4 ��eH��:���X������U�`��yߧX:�z���z��]X�ą=�� vz�N4�Ct��Z`�S�n���-���fi�w�+�|E�Uc<W�kÃ�ݡ��N��[�%�$�=���e�1�����D�c@
��ܣ z��V�R����o����t���n.�V|A�!��7���#�[ǜ����f�#��Nl�1�e;ô�[�sdGڇ���ds����n7�=����w'�s[��Ɵb�+�������,eoK���'�����$�ݙ@T���U|�
�&^�UG%�L�2>�/9�Ak�Ī�%��A�<6Eei99g�pz��hǶ<��'��D�˻���e߽�\�� h`�b��~��w�2G~��gRՒk|��"߽��p ��CL�o����ɏ�$�b��g��·����m�C���"a��u!��}{�13|(�V��w�����Y��'�g>����Wy6,��1��h<�v;��4�+�1�ˀ��>��1Lp�C�*T��[+��Є���l�F�3�3��Wrf��M0��(�<��{UWg�<T����kFw�c���ġ9�z�V#f�G�8��bF��*�{ ?pzC�9|�QJ�`A_P�9n�!���k8�\�RX1�Ӌg�4co8'��8տH/���.��ocF��˶����@2�<ώ�1�oE���{�����Y�c�]�.���R�� �R#�W��;�{�T��e	^�ţ�, d�HMG�!�Z�+ه�P�m׶����-]vC(/�oy��J��L»�0�� ��(Q�"� 8��$g��
4^��i�d`傩�eP���r&�M�U6h�3.���� [X#O�qf�Z|�m˕���W�=��
��c�Wv��|M�ݺ��d�8I�*�R��=�@����^_��%N ��9��KݴX�;w��f譎N�>O�tBx�+�����.�̿.#�udK�y��g�7�w��@�h�sZ��Кe�]�}��rt�(0��8����7�K��V#�Y���1��bV��%�d+�LW�6u�q�Y��f	|������M��u�I��Y��6�� uYM�8�^�R�y�j��%C�y�rw%jSx�D���Յ�����O��h�7�4I�l�!�֪q����t�����&���E�ZNB5�$����x3���d�ǝ�u����HS�n����0�%)���[��63��y��_:x�X`ѕ?/Y֢o�[-�d~h�Q|��9%<��3p�ˋ�/�i�"��?pv#�֊=]��e���m����ߴ+����L,��b��4ڈ&���t$��;��@�u%�j-p�ǁ`��1���J��h۾���Б��L)��v�I�w��Zp]e�e,W5EC�/��k{!�F�̡�0��a*��8i3�qLN�<"=��1�5Eۂ�7��
�c�7wS�`!������f1��_f�,�>�`�p�?�)s��fI��?�����=��%r�('<E���py�YA5Rͤjt�����^d�|8������ �0��4�Sk�=b�<�C�u�%��gۘ�:8!��K��>���^IA4;����ew�12���\��>y��^P�:i+mμzU$�ЦI����S����.��y*��\��m����9�ѽ����B&���~~��k��)|��i���]���2Y�0pbk�=O��Y��.:Ai�j�}~�t���.�pv�ߩyb���Zo� D�O�_,xͺ�������r:}�z5�LY�!�!�@��H&�ɘ��XU�Z��Yt\��͟3���;Y�<���}d$�Z�a���6k#���K�Q�ȃ&�?bIzt'&���<�%�uyD�V��Dj	'W� ���P�mt�����3m���~��tkAZ�4_�-��6��%d�0��S�J�\��L�'a$��77�Gt�O"���u��.��^�"A%�(�4��[�M(�:��%퐣2�p,�G�B:�8"K�3R��ŧ�Z��I�_��4+�.��j���x#3 JL�7;���t�F`_��l��Y��G�I^�hp/�K��!ۉ&��u���\�Y����]�8|(8^RpƱ�7WD��&yk�����i~����̀�8�q>~�p���)S=�$A����P|��{�����3���wZ�=&Y�.48%�ckX	���	GX��H�~2�5��������=8��8� ��M�l��'�tu��~�̞L��9 ؽ5�H��5�Pa���ܩ:�׿A�Sc>�x��t�{6�$%��0�1��d���9��>��p8����� �;P�Qz�c�]Q�{�@�8s�Pͫb+�Qͤ�J��%6��@�u�ղл:�YGr��l��հ�c����0(kM{pf��"��+C2=�o_I$e�|U��(w���o��+s4}j%8~�z�\��9zE�8�Rz%*�X��(��F�A4Zka[�a��{,���Z�YRa�����jeƫ�3k}��\u�Ih�.د���.{���S�B�����c��8Q����..��<rV�rw� �op5�4r	�Z1�E��:�M�o75:\h���9V��L��"�k���C9����v��=̑�O�`+����@��X)
T]��Dz��=�IH]ٝq��s���ʞ7�d��|���J�\�v��=-wUj�~eQ*������=ŌHC����o�"��5Xh�n- 3�^�(Ŷ�� ���UB�Z��a��.ם�)�U�t�G��@P.�iU?�qL����N����r��"�:�^s������I���~����ѸV���҅�8��V'\�F�\�B-�3��T���F�R!�D�V͆��$~V���ك�_�t ��B���~֬0��#_d�C��h�@���FՐ^����l���3A��A�7L$�5�<`~m�Υ@�Ӑ܄pU�����:�E�\D�F|h����4�ڧ&f��WE0�"�ݍ���bouu����I�`�j���7Վ�#�F�	���w�1��wEk��@�� ����	�+4�V�ΞF�� �c �w)���F�N\�����<���ب8����na�0ހf�)z�G/�Q���H����Z����M�P���� �t��;4 l�E,�����^7���*!�Mk���l�_�_��,�dN�/۝���G�l>�J4���v�}bN~�b�:\� $5�r�-^��օÞ�r��[���uW���2�
bc�R ]oFX����g�/������^SA�[Lp��K"��! z}5@/`��ʢa�0U"�`��T�v���S_-U��a�T�p�`�p��
;qm�m�]L
��l<�a�bH�{~j������%ُ�8���S���VR�]��:Շ]pg�9Kſ/��aH@ޖ8|q�Ù�AAJ?h8<����9	"��j?0��,�A�c���;��yp�.���-$���׵�%t�W�)��1�d����u1�qh��Q�,<Nw���`��4�W�>��KD�,H �da�"L��������(Δ�^2�
�h��DJ��jn�B�w�����qߝ-��oc0�t��k�n#�c1�7����4�R�E�[K�Z'tV�RX�/�Ŀ��U�����gӫ�x���뱪)m��
'���H�͂����&x���������lo��v�������B�;!
[0��.G��Xl���w�T���	Sq�Vv�h���K�� L%�>�g�6;��{�T!WG-@�bY���,�~]�����Xv�3�Z'�iz;���~L���ʷ���3��>�pe�+:�{���N�'Ȍ�["TEۡf�%Q^�q=�&���/�F�3�Q�dwn�*kK��(�KzW�G��|���K�d�Cl;ZR�KOi{�J�L�G���]XE��z�ܳ"~R�+�l]B�Xh��30�Kq}cTm�X֙�}�Hd��mMqa�'�tCa8e ǰ=��~�x~�n��U�%��:�nsp���P>����տ���5,�Н�M�\e;��s�(P'���ֶ����j�&0�(��D�]B�$~kzeu��m*{��;�w�ms��c���H�Q
X�⏿�V�u��\j����(N�b�1��+�?��g���yǚ?c�څ��[�ҭ�T.AR���`���ˠ�\���+mFT��T��������b��0�������5�nTYRn�<u	I��"q��C�o%����T{�-նo?�HZ������酳jo�a�08���z"0ǭ��S�N\#�N��Z�qF��V��e��y�6'*�xY�50}qxƠٿ�P"S	��1L��@�Px	�h����Ϋ�V�')�7^.5-s@w���ɁLs�a��3�jUġ7H#;�4�
�i�<�tB࿥�����U5i���[��$�X�t���Yj6��Tsܬ'�
����!������d�����פ�Vh4*�Q�~���y���^~�t�<��-�I����ߎ�p	Z�浴�K��خ�d��t��US8(�`�_R*�J��Y�L�V��z�n�u�WsJ�dU?Ĳ͛I$p��"��)mE����	4�	V{ԁ��N�\R���Y&u�����(�~�\~� �5���bA����Ջ�@<j�.�rZeZ
����7���#I���hO��]����(���� Z��x�CԱmHl�'�hS�M`+kN��Ͽ �����'>桫�r*��D���OG!3��wޯ|<�Q:�n�^xգ/�r��|�,�*ǀ�c/s�_d����h���y(�Y�4/W�SS&���geD?��.�i�j�9�B0҇�g�s�H2�˭D"��[���?����8J�Ӛba�!م!D�r��7��]�r�P�q������k�g�ݟY�2/�4(RA��� )ɡ�2��}�U�~�����E�s�6{�?jɕN�1�?ҝ�^�&l�H@�Ѫ���{�x���q�Rģ)� �v��@�݀X�~�+c��A��A�H�"��a��aYV{�B����Q�g`[.�;�p+̻�~�=���E:-�ъ�Yq�%��Z�i���&���k�`��L�K���J�ELH�7X�!b�����(T�G��>������?��+4�(W?h��aN4jD.��*\����1\n.qR�$�EŎ\�`���UN��K�Bw^�%D�%�^���i�qH:���>:���{��"��J��0&'���Ʊ�� �����ah��CƗh߂4��'%�_�ϫ���������f�N����r)�(��<u��f��t�1=��c�æ�.ä�ya�{7g����$�v���e�G�+K�u%[�bt�n=�N{�6̨٠>Uh��J�hn`;P�%?L��,����YFew��e]�G�R��Ϣ{�5��cK�v�c~�\�5B�G�����M�m#I�����Q<DO�E�jJ_E-b�Qf#!U9�f8,DM�Ll�M��p�Bb���,+�[��T*� �X�������9:��N�)��*�c�w4��a,�=K�������肙��--%��ô�,�&@����F2|W@��6=b�>��������k�B)ս�+�CD.���u?�/��x�8_��?��&cw�I�8�6��B�9'��i{cE�o(��@(���������(4tf�Z��H,�V�SQ�Q�B����p4�����;A
�+�@�c����:��p������٧�	�t�ǫ��oVyJ<�a��5T��UF|���T%���� j��&/���u�Eyf��n�'��Ǉ�"�������`τ�H߈k}TW� �R��ǥi�2���wN�D.�^1�+.,0�	b14�u�3�Uχ��*�����`f����A2���'�FD��Jb1P08e�8w�gEW��������|2�){�3��y�&�̗�s�'^�DM|�Ȃ����v�D�U������vM.E[]V�#���.�,u&�KCM�E���y�3Bi[HHi�Uwj�҆�p�s�f��[��!pB�-�Ϭ�){��p'�I�礄<����m�!$i��75-+r�A�R�N����x-��gz�#Xt�:��K�bL������ר|�8�Cb��.���떢�ee8p����v��%q�^D�Wz`��s�"�
&��C6�*#/7�λ޺};�[���Y�����
��Pb'�T����X���l��&����ݶ�����'��x��R�Ê�=ՈM��Qs�FǞAp&'�RNA�*���m�=41���	�^P�4j�
�x5�>���~Z1���v�7���=t)����>�U�b6�H���w�>�������εV�5uxO g��"Ӹc&2�2SU�z�� 0��v��0��)��Ze9�k2��T�˛L�g 3� �o�x^7I�;Վx�,3X	9�-z��5��� YC*e���������G�<�>4���&�ϖ.�U���|����?���mŦ�<��/�z�Y]�Yti,%���]�����js�!�Yu�'�͇��ڄ��}�^7���x��5�R߱�?��=U�����Z�Q2��z�,�	��:�*=nmП�$�3?�<E��Y4%�訁�_/��t���#wL�o��ך��''��ڒ��cXh�UOh��FP����{�U���]Z�B&c���i���f�0�5�r�(*����<�V"��a,��MZg��*��EF�K��f.����97�=�~pN��=^܉���$ȭɂ����b��-)��4}4�R:���PZ�C���|���ZPX����q]�=��߮�8*�O�Z��[��(6�f);��P(����h@�ߍR����Cߎ�K]%���RP���@e�5��Iu�,/Һ�uϐip�%3������qJ&���dpNrn�9P����#֗��I�>�
�'��T�l��,C��I�"W�%�9��ݠ�+��~0��垼���:�����E��A�� v���<3�u��H2Q!�nl���-S�d���f?���݃|��Ѹ
H�&�m�wlL���ͣ�ghHi����/�K�����çM����ҥ�O�x�+��
��p���<����F_I�q��� ��Xڑ��)�.Iy���,�O�;��uA/�a;�!ڛa�,
*�3П��bG���0-^���=2y�n�0�bmR��a����ԙ�o��_�Z
��?Y���i2x������ 0Ih;�����!�$M�7O�gh=/��/��E,��b��L�/Q�`&b'���]#��u����)��7�C�K
)�v����&�PED��_4ӻBx�?���?�>���"���۞��v���~``s?�$m^�c���(8�'x�t�pӎ��م�P� |�-7yZ݌���B���II��j��SL�9��ϱ��a*�CH3u<��^`�8��Et:ǒ��2�5�����DV',��D�)��F�N?;���e�P�;��в��Q>`���i~ Nq'�]T�XJ�6[���+]*\����]m�W׶H
^<�������d������ /�pq� \��h���feR^�����f��K��������l�k�Δ�:�a)v��J8c ��ƞt�Ѿt���@���Rfogu?���*�h)͸���؆�sm���3�v�b�P���܀�s�x3wJ���4�����o��C6��i�T%�T4PPT�(���!�M]_�ajO�\#�R��p-��d^�8Űٟ/�\ �J�g4d�f�?sFg�������fuIiȺ��o�/T��&�-�a���ː����Ǵ~��(��L�P����X�-3���{P�+���d�6��D�������������n5g���zE��Eѽ��{�|�����L��:u����oͨ�Q%�B�V�?97�T�V������ex�_S���E��S@O�5�:8t>۶Zb�˰&KO�LA�T�YRt/�9��~#ap�cgoAjX�$ߢ���Br��:�����h��3������<�����g烵�M�T��a����s�Q���;�W�zs�vy
��:�\I���c�T���ֈ�ۨ�"�j���qkob����2��]�����gm������G�VS�o,t���-;�-af��`�伧}��OR���'�x9�3��'Ј2���i�R��/��e�|�X�,˫3 ʬl8�绬��c'�,m
]k��`���t�G^�"{R��i��O��3��Y߫e�t�O^\z?�i��(��s9l���c�0P���޴�	����U� 9��vH���$L��:&5�.Q�!����`��Ή�/�)�:�t�D��L�)�
��Q)�U:N���"��C�j�o����C���R���O��?2����o��U�,|��(H����#Ń�>��� ��'CӼ����1W%�4+�Ԭ\�b
�P�{�>< �I�R��{�x�Ėd?Sv`��^��RɇȨ�M�̹�� ��2���Y:u'��c�Oe�y��ck�>�BI��>�s	�/�C�%��ڞ���/�c΄�>��,��?�ˈ���T��F���8������O���$��/R]�֩�:WǺg�� �Ƃ}�D����J;�v����EصP�4<Kx+�[�U$���>\x�������MI��`�)��b�ă��%^G��p��'j��
L���O8��E6)˟�Ѕ�V�����D��܊72�<�VDG˷�\Wsfjmf؍fd�r�L�P��iI��^C[��4�U��*�w3$cL���2�H$���7A��v�Qq*����4��ǲ�]:��x�h��G��? �E,��N���t4���P�ȿn<�g��(tc���ވ������#_D���5D0,b��U�4Tzgi�ǻ�7��aI�7�s[>0CM�ƦXkțp��I;j��m�47;���2
���QD8�h �|���}�����ہ7�~�Fc'�*T.��ע��s�0��J�F.P�4Phy�{ŵb�S��Q~h-1wM�A�aq̐����X�I���r�0�O�T��Rsg�G<E���������!Uk���I������#�?��4A��8�^9Fa�Pp��^�(էӇ"���=�W��Y�L*�k�p��7�h�
����Й�:8s��dY|E�a�i��1&��,р5�hH�"ĉp�"�b�����;�l&"Dtb��o�kJ�k�Iq3`�II<K^i�q�,�G��1�w�q�U�V7/dk,:��j?hj���r'�L����N��!�2���5)��m^��(|UG���l@����9���������x���#S������2w�lv p<�8����'����o6��u|��Ee�L�դ!�hsh�M��h2��UU�p\
�5.��,��e��$��ٻ�� ol��z�Kk�8!ps����:+�&$#�1��Qi�'�"/�vc�ά̀d���v��-�MdhB���~���7u^��9]�h��I����u���/Β>/$<�[�Ўh����i ��Q{�B�a�ؒa~�?`o�.D�̫j��]Nr����"��E;�Qx��Ԓ1ЌA|��X��qPٷˊCL�ˬ�蓦��=y	EV��J��w�yU&�-�ǖ2���I�0o��x|`�
���k�.�˺ck���&�s+���1fW��Edt�(�J�Dm�'!:�p���c�����l[�2]�M�=b��x�Xiz*/�է�ư�"��G_.�h ��\����D�oX��N�DRhϙ�޳3�0��4o� �^7j�̴��u�~�n�/��M�����x3��VQ`]����aztK���U��Zh�6A�_���
��;Jg��C�Ց�PrWÓKc�협1�9�ƻhr��U��]f�Y�ן���cj�Ư}H�ʲ�A "]VM�4�'A�CJ�;�A��x7~�K�Ͷ�)i�����n�[�{1��#���r�ʖ��q��d�?DT]q�Y� �0�d�Q�_`�.��?(^�:@�F�L��20���dR�|� �z�1��4ns����+D�q��mA���E�4��4��`���Ch@�1| ��	�g��"ێ�ox]M����$Y ��Q��mz��
�o ġ�0b���Y�ٓ%)�/;� �+��'�֮�Ⱥ��u����
�銷MU�E2�K�w9���X�;������$	�!��P*Cv-���%v��8�U1��Wr�ȪRF^��|=�;��^ÅSAˍ*�Ʒd�SH٤�@�Qr�+�E*u,3&J$҂}�6(�z8��h�-������o�*x���r��jJ�i�����Q��F�䝤Uq�bzҶ�*�Ѩ���
${Ϥ~dIW�j��򂪸�R� �~Y��-�/?�u���#�-��7 �<
�s�YG�D�1o�4���������KC�0?�Z}r�҄��l���*z�! �Bg���3�spZ���)�������"dZݳ�����Y�)�ȃ��p�ѐ��h&�?0v~����l|�B���zf
����w����ov�'�}���T}����mkoa�"~��[��������s�,z���`�c)НLO���@O��.���8����J��K���4c9�{�]�*H*���r��Rwn�c��kT��b�cT�!3�Z/�D�Dl���܄i�<�Zc�ȑ����0����JX���� �,��G�k���ǧ�@u��m�`]��ùT���Y&zf5��"{߅w�j���V�0/;C^bݡ�K��o�V�B��M��m�o��l%G��za�Ė�����	�}hB��3�}2�4�d��e��qB�>�����.m���Z�_��xny�n�آ�Q����B�	�M9`v*���"!�h������芥/���}��7�k�T&���`��-��YL���1�@�{R���+�M�Hn1� y�M	#p8�Kwp��+NPU:�>]�����ɂ�=d��o6�Q�Z�����|�S�n
����}�0�h��->���d1�����^����w_�݊ʩ��[�<�u$��2�;,f�Jϵ�x�:�c+��$�/!�|�"�I=�A�m�7K�# �P|H�o8IXw�a���('⋥���1�����pӌF�
�����/��ҿ4�y����I�G�e�.`& %���@��6|����Q�[2�S����,M���;EO.���~�,����枩h=�E�����Y���sUB�7|�i��bcs�Ȅ�Q� M���-1�\�EE�}8:��0��[��آ�v��0骘�OYU�� IV)9e3QXl{�e3�yEa��	�X���)��c���aB�1���PT� �����}�����.��`a���d�9:dw(��N�)X��O���/}+b�����2m0�|Wƹ�+(�U
h�@&H��h�"��6�a�c��;e.-.-߫^
�t~��ܰ��4��^8�VH��w���<����6	$���ז�O�#�>TRF�~�r�}9e8?Kν-�q��c��a��e�%�ܹQ�%O˻Rd��)\,�~� =�|�A�˥/�������W����Ԕ���=(V�xq�(�Uk�]��X*�)����Hp�z& �g���@~M}\��l��/�\����ڢ�	,�R6z�ӺW�]X� :}�؇��f� {܈ ;?�����1Y�q�MA�ݮ�� � ����:���
v�mk��oү��1�<{��
�#�����ZM��v;W��}
ZR��ݶ�E,YR���~���HDU�{礏+>a��Gh��J�W@j=`x�����zS`;�p��`����q���)Y�q3�)Y��]�ƌ+@sQL�M,������BQ��?�9,�\���z�9z)��ŅQ��CLl<R��6B	tH�M��:ͽ��r��_�7�{�8�?�e���%:����¨bhI���@.�>R���c�x�d�!&:Ԗ
���}j�z��˒��Ŗg�C�R��6ѽ��b���1	���şC�ǌd�}��+%���I;3`&�l�������8@|WG����#�)�n���	Lj~^��'�kxR�"�'�n���I��-"<���.����<=m�c~��Ɉ2��[�i
��f(�bp�`V,-���#���ߠ�* BM|���JC���7w��t�5n��C�oP�x�����kw������'�t�NO���ӗ�=�}��H��m��_�1���a��Ɛ4mK#��]hU|*�����w�ê�:����f�>g/�9�ǭ��|�]�OI�K!D�У�ػVW��v��<ȟ7�/{fA����B�ɏQUЖ���~<�<w��TE��?�M<jj�6���~�Gq#p�����[�|�OҺ#6m8�-���:�h��L=�U��"M�W�����̨Q�L��_����w�m�r��cr��9�q�􊅝Y���{�\�m���qF�깱��W�Ib�*l����9i��
Mr���%i�9�NL�FRF��i�e6�Ϲ����s�r�~j)��28��8 �_�q9��	(�*H���r�^;�|�0,�WCs��";������k9�膪>�*�Y�R�=^��Zȝ���5�:�i������/o�?4E��0��[ua��:�������AJ�	�#�(jJ��/?4��s��P���>���5��"�)�o���h���UG�4TH�ޞ��3w���I�"�k��pj���㘈̈�jOjF�>+�9�Ն���Eآ
�z[����ƅo�]U�R��c��*T���O<�)["!l�l��K��YK��d�햐#�\�#��3�o�U� �V�~i]k�⾽�.r+�Y�.��F�KY�'�,Z`��} �̷1��D�Fx��i�r�ƴ`�ozFͽpE�n~�ҁt?6�ֱ̣)����(ً矰P�Y�.���wv��
'�b\X�y����Ç�F[c����E�ެ4�Q����t�"��YT�Mw����~&g�1ì�/��a�j0-\v]���[d/�0@�Ґj����ܿ�okK(��'�����S)$s	[@o�HDb�eS�vf������Z�Y�Y�bSů���qy��L���5	����8�ij>+ؾ���	��,���կ8����{Z��m����PpGl]�uDĤɛ?�@_���%���C�~ըK�x>/�.��xG�i��R8EO��uh�@�Ů �ɅL��m�$+���*��M.�VH�$\ ��"*�!�����z<�_�Ҷ?kR����̘���e�&���(`���F���1,�m�v���u/%��	�q�ֲ��:��ڣĥvPS|�U��� 8�_��]������@?ʴ/�;flh�i�Bq.��dM�L����l��IWa)��u�km2e�V�U��Q8��f�����{�"�	ف����L³�W<±�v��m��@����H!�Cz㕮&ٞ��;�XU+ѩ�f��`��ze�#Z_hZ�Rh�����W�T�	Bzv�L"�!�%�@��o�M�'E�t3'h<� ���1�$������Ja���+(ݙ�*���_9!�h���6`0���}���N,�����|*�͢���=k��V��Jį�3�P�G���C�g!�5+~�ux���������̐|
�L�j	Yu�
�D���dǌ��[�̌"���Xy���Z$-���O�5�� _#�}�I�}�:���o�"��vHq��Uʜ 6�	h�Gj��1����j��i~���ZR�k�����r��ς"$/�a	eۼ��&r�������?UT����`�c(��=GJ�2�$��������������	J��gw��m^�āDU���jD�&Y� -��
z9-?&�:���Ԏv����Rc����S�p�c��_+�% 7M�Az�D0�^Wf��W���]r$�}�~�M��3̖*��P�X�D8�`��@��QD:&�{j�lK����1�\��h�$���Z9��qU>�_r��\�0#�m��(
}�h�Sn5rˋ��Z��S��e�̞�3�P^4)���ϸ��/���%�����%��J>P��@�)�(� �7�ͪ:�oe�ݻ.Lu�x�B��{��Y��F��^f�B�? ���'tv[����b2�����_��b���-C`0�ݼ<��P�(��g�^���8Y�[��L�t"h�/���\��k����]��޽m:T�vN`�������z�Zw�J�Y��UNs��E�"��;�h���8��W?�-P�=��A����_LTp��EDyU��j`D;gi���r>������hb
�K�L�ċޠw9zs�b��zʅ�A¸%ܹ��<&����R�.��e�!�)��Z��s�¬P���l=C9~�aa�|x$�	�P��p+�O�o���K��5-�>L�ySW������8#����t+̵���7��-�7�P��:i�!ՁB`�VI�S��U�jy�\i�sM Z�"鲩˞��T�^�l\nze�\Y
��T��ph�����-�ț�����p)&����C�E��|��	���;Ӆ�$9&;k7[@�5�ȥ1��y6U?B����֣�5@֋2�D�gIQ��D����+��Hk�j7��!���x+	�B�Ƴ���V��wP���n�x�>�v�S�~�b���u[Ɏ��H�:B�#K
�a�2��Gq3-Uzg[�}�������gwd�/ܹ�Dg�]釞$ޒ�szP�;�}g��� gKO�K���F��EP�� ZH��Y�}���8�j)�#MH��׫��pS/�!�� �A�w;��� �X�S0��D��/��G���� ����S���@ �����){�ecʜizR�x6ʕst���r35?�av�(���D9���g����˪�����xg��X��|yz˦J��>(O�Yz �F�I)��N��nk����;,�]��l5 !�����!m����� #�����o�������^�k�/C�S�$9���<��@���J�q	�����*:ҍ m���
��6�-P����n4(��q3*�X�x��X:si4D���L/M\�1� k�g�ؕ�$�� Y%)Kk�9��԰
_�-uV�\!9�"�֤}�I#���b��J���>��YqAn"$�u@��������\�m��O�!m.n!Dv<S�:��"O�\̒][<&�g���@���y��XLߎ�] ��Y��\7q�8��x.p�C���y29���2t����O��Lj%��b^�!��5�ؽ1U	В����54��|׈��X/=��O9��~WR�,���w�AP�������8�Z K״ys*���&Pc�j �&�cT,Y8�ց�|ZVP&��m�s�>5Y�;t��^��AK[�L�k���1T�E����=e�{��Օ?��}��Beق�"	�ƙ�9^�Z�\H�2pI1��?>����C�*a��|�Q�i��S�P}������ �^���Qa���-i���вy�E9ؒk��_)��s$Fy>�?ɼO[ێ4�[�Lq�{�e���6<`���B[�"ɪ {�ms��q߀��}����n4�^���kF<i���.e�Ut��d;�&|ڍK�v��B���-�H{�PD�a����<X4r��H�+
�^�l�5�#߭s1z@���↹�,7��u���G���Vc������uk�j��R3�g�l]墬>���X�BC�U�3qg���ۥ'���� %��԰����n2c�5O��h9!�\C6���Ŷ՘Rt �m�ZȈ�eX��ɏ�=�b�ǚX
�:����K\���E���/)-�����۠j��s'�=aE�F��z?y��6��櫀]_A*���&�)9�h}��^���V=6C�L؃	�-M��lT=����M��	�w�|�%�$�)�g>=</��C��#�����{8:�*I̕���K O��!]�N�'���G��j9k�^��w���C�pHo]��d�v]�,��y�M��Xx$�/~^o�r5���Lb�c�zAA�G��K�J����iC.��3Y3���"�9��U#4���_,��Ma�.�doVBAiy�*���G�3:9�!o��$���s���)�F��l/
�j�բ�۽Y�ok����$U0&�W��9�+�X�i3��T���T�V@rMT gm�O0���s�ᠯ	��8��Yr4�@�C�$�/������r(F��Y:u��}e�%WH����m`�I|:��r]t�����݋�:��f��	�H��L*r_5��2#]&'�_��&����T�[�'^�����z ���e�L�O�9�Y�T�	�J6"�Ǐ��>�u���TM_{(��g�e�u}��&8�4kD�4C��{����A�6���.�v�q�	���9W���d���.��ڡШn⭀-Ohy|М�T9�v�nQm��I����	w���.���D��r�@Ƅ�N����@����$݇��.�3��+�A�5 XŚ����O�ok,�?u��7A�;^,̈S�7��i���r����":��[�u ��x��G��h�c-i�rS#3 ~����i0Q�`�G3�io*N��Xf�e4�x�b%Թ�D��2�:M:� �Mjt{0����T�O�4?9����-T��������bq]z@�KeLŘAw?��hh���B��j	� v��U�4c9�>Q��qu�k�2��b>��U�K)s�0�]+�P��Q���C���-���H��/��I.YI038�B9(r'r�y��������V�1#���UBgс��辇B�F�XI0�m5�E������yt�"���PqN+�aK+"��R���N���Đs,���	���QЁf@���W��|�I �{����)[�،җ\#������Hw������a�'+wY��˸T55kl��0���1q}��Aa�+h�{�k:��u+�� 1�05�_*������L�E.����ŋ��F�H�W�ŏr;�3�E =�¡zEL>���龜� ��dܦr�T�hO������Z�*�`��P�H�y$�$�n���]�bM^Fz�gDf<�y�GA���T|�j�l�,оմ���[	�(�E��kEz���(%4!��J0��Cx
��lt@��:h��@�)a�Q[72k���XL�.�O��^Dy�2X�' �8�(���@�Dw�-�w�?����&��9y)S5(��B^ $N�N���M2����{�س*�\��,�u!�d^��^�����V��K\��%z�u�"���I�6<3BB��m���U4�0*�̛������$�z�W~&{����Zu2�����Su��d/��J[�D�@F�}u��`x�U�t��$1/�Z�l�l3V�#��Z�ߓ
��ɢ�eSDoeu8�T0w�	��q3���ǔV;=P��7y���=�!+SI��-���BW��4�9�NjJ4�i��ƣ�v��R��[Rl���eH��@�a����՘tES}�/eV<#�@�8*D���QB����;?�,�RP��n����0p�̾�������H!� (5p��0ܒo|�@�Gw!d�O6���z�0�<-\�Xr�s�
� ���$9��RD���w*'��B��4�����&Z���c�mC"k jl���+>wP)p����X_
�4i�Q�:ܕ��^t�ټD5��Z��h�&�Oc`u���ƕ�{�V�v��kW�3�]�*��s��^���0��A�[D= e�ΟJ`��;���S,���5�E����w�m5��~3F���d,-�]�"��	 DN�b�w� "�E�V�������,zA��<U��\����S����u�gק���K�LQ���1ȉρi�4{٪��L��<K�%���|�4�0/�<�K��x��.%������FP79���{���L�m�.n�S))��S�g�W���l�C�_����R/����.�`
��SiU1p�&v
v`��rX��"�q� ���`����@�	2nW��8��5����K���3&��=]8b�(K����޻J��l���eq���J{��U�~3M�g,��k�=�����\�Xq�8([�U�n��/n��Px=VPY�����O���oiw>����`R��rä���iFX{J��)"�
14�y��M � s�'�
��������RT��V�;��Y��[��A�vJ����fY�L��ڳ�؃H��RW�8�/h�R�ur܀e
DE�����X�]E%)JmS��"��%H�R$�id����*
����w	���ե�Mu`�w]n�q2�b���������T)z���_]� N씿�4��>�{��	]%��#���H�0=x���[�싽䜲I����$�ݪk�0x|ı�<C�����h���Z� ����*��#`e��}� t�X�x@1���cV�}�=����d3K�0_N*gK�����f��A_�UY�Og%�B6�H(n��2[ 5Z�s��>V}�*-\<2���}�'�!�W��
�mWc�sR˛��=�K�a���E�i���*���1�c=W��2L\��~��B�]�d�\b��z�������!b\�l@=�@D�t	�q�R^��������� ͺIP��;�zM%2+͊��Y��W���c�
#ߚ� �8��\Jc���]N0s�vK��'�A�%��9��;P�;��N n��1��A�.�����o����$:)�Nn����=�'�o.d+�s������X������� ��ȹ��S7�����U����^�>l�bu%T��7�c^^���ۖ��g��΢냶ܾ~ ��J�9����(�� �q����n��{%��I,x�Q2<�J[���I�$����ɯ���z�PPje�?q%:nK���I����%�;�y�|WU�����o��_�N�پ})�&w�;��&��0Ջ�݆�3�w�K��*�������şH����4��T`ἲrH�BptxAփH�C�嗃,���ɮG��#'(�McP��Md6��a�����F��c{���8y���ktwy�� ��&:Y��Tdf�?�G�|`z1��X�eL�:U�G&�3)�G����"Sͱz,d�RD�4��
��z���#���y<�	���Fr�Q����a!J1�Y����ܓ��M,eD�H������2�Q�Df��ӣ����~ˠ�UCF
',]�7��M�ݸ�b�
j�Ř�`�Ꙅ�gQ8�C΢8DFKmƳ+	أ��!#1��Ѽ�e�B8��Q�q��Fsho�sl�A�G@jA�  �fJɭ~f�m��o��ܲD!F�mm��kg���Y}d8�5�kF���B�p�o�$Nv�w�O5��_ �/��A�кTS[|>9k;2�Z���f�qt`���c��`k��S,�������s�5U�@�{;�=Cl\S�̹�W�IHūj�Йc����\p��t�ѣ<�a�J�x���!����'�f�O��n2R2S��u�ux�j?����R;0S��B����V���U��MH�,ֶ�
����6�� /��ǆ��P�GA�R�#0����7깃f�i�wo��(Q}ƽйMː�k�zCz�<虏����Dc�}�R&1����k����Z��.�m���?C@q��p�����a����vH��3qz��ذ7CSݾU���@���R��l��p�~�$���*X��8�
Q�ࠛ����y�F\�x�ڣ�A�*}��29sD�'��ExVi�c�4��D�u�E��K�&v�@�Yќe��>��,�Y�[�L� �⇧��A��.�ºm5 3z��g��w����zR� ��i�-��X��^j�߁4�H��@4�g�9��u{�3�_�[�^kd�1m�l�iDO��fA\S}A0��<����
[�tT������L"b��0E����1�#Ƌ�Kug�t�n�Zg7,e�2_O�+y.�9���)	V����D\EB�G�h��S
x�M��Xt2<�����iֲ\r\N��n���"�T��7Ў6��	��
S�7��t扈8UU�٦����>폎��+�k ��_+zx�f���91�t�T�쵚'b ���$�o�_���Eq�� 0��_�F����:%S�9t���
�{E"�uhr?�n����~�֮$�v����X'��pY׭�F�u f}��$q�r�7A���Yn8(x���H@~��Z6��{�������@�yZ�3G�^�{�t�zb2e�Z���|z{ͮ��� �h���ԑ
�MU����|����'�)G� �{a�)�VSC����Ǐ'�D��^��G��u��
��hR!�vL5�UDdPE�� m�C�LJVVbR3&�9�¹�l���bZ�|8R�����(����,?\�q{�P�' � � �%���ņ�;�x���j_(�y|��T��cB���#���gF�BgY�y@�1��������Zi�l��������H_~'-�j�v<�(�����еB�mڟ�����	V����Ӗ�a�{z�U��~?��/��1�4~>*V�`x�0�L��#��Y8����㇘�Q��[��n����Z��۱Y'2��e�\�2�ҷ(f����I9����(^��n�K������/_�
��wK�Frd�4���&VA�@!B�w0=�=�'|U���wfN���=��Yj��'U��]��I�iq�
�{L=#sSl_$HŌgPB_����O�?%LG������H���������"�<͙�2�t��IvQ�Æ�hK�aV��őGP��2��:����Y��}(�$,l��"� 3̮�/��T���\�Rw�\	Yc�o�B���b���5�;{9�TloB��S�+��f��	,"ʍ�I�0gw��Ӥ�'��,��� `�t��yǖ�l%׋�_|�3��n/�G�uGz^��w�y�a������<5��'���
)�s��b楜̫��py���p��j����{W�G¤Y���p^�=��,e"���K��h�M��z�c�}��m?|�(��ٍ�8k�ᒼN[�c�$���Yց[��s#}PN��keb�Z��E<�Z@1=8�7��i_�y���p,��ܰo��۬с ���4��[SY-B�.��N�,�}�V�6�?;2r:�PPH�y���D���S&8\�7GPZ~��{z#��G��z�G��e���|�2��+p��Y�?����j����6N�M���>ʡ5 %u��ʕ8��Kxͻ�W����wl�+eD�}w��W��Z�*9���>�v��� ��l�w�"5E;R-8�_�{J��GmX'H�Іט{S�ڛ����LC`�h)7	��x�3a�ꖄ�v�Xv#�
& ��{S#�/R16��X9e��ϲ��t��^}���t{�T��<��Ҹ�LHt*��d�DkG�tz�E��-��fq>Sp$$_�{{��ߛ�nC%���e>�*��,��B*��؄Iš;`�����_�ϋ�b�����σ_a[F�BW���D�O ����pF�.՚���(���zլ�k�k�3W^�)�~��j^�H�*{U�m���/��K���nt�����n�<RK����������q�,0�zi��1�O��Zu����vEc�����?���ğ�&���3��>;��� *b�yI�ʑ9�	��Ov��KR��\��EM������� ����q�7uv�����_�ݐ[1�8��צi����I-p�0����q��e}˱����oq�NO�kxq`*�D���,�����Y��eǇ�������!Tb���ڜ���՟�5��B��'ġ�U��2wskh��YN^�I�
���Am#�u�|��;�\l�wZ=�2"��7kܧ_�ޘ���.ڑp�w��Uq?����֚��Q��G��t�
�s����䏴N����9� � / ^��(���8q-�i���c�v��@!I 5������kQZR��ݥ,��フh�˹�K�j`K��p�c[��m� �6���uH3K�����{��o^M��qZ�����,<˾~��p�U�y�wԚ(6�`��;�er�s�9
���+:7V�P	H�<M�Rt9�n��W`ܚ�6"��G鶒�2�����7N4��b+��0>��rН��կ���^�)�J���b��H���s/�"��!��5o��:Zuԧ��G4�~7��ucI�m�i�\��n{<[�!詹�ޜ�1Cg�,Y�����Ѵ���d����X9.t�TYB&����f2���d�߸���Z�Uz�k��'�$
ҿW̟/���5X���Ѿj'<?�����*�m���9�H�K�٤'��}��de�<,�j�{O5d��-p��'�y��ĔF��	� O��n��x9��n{�T�`�I�=<k���GZ��R�I�&�޼�
[��9� ����#D�Ua�[`��ܿ��뢡 e���&��%D�Mo5�mF�Zg��gAl�R��܌z��=�8�f.�xS�R�Q���m�)-ځ&x���9��J{�m4}�=�#��N#��;ʽBAa#ٵ� �֑��P�^<3�#�Ae����0�_�~���ryc������#�i6�=R��J�Kji��l��$|G@-'���g��eߒ43�կ+��d����A\ȱj�J	�aJ�ey�^TbJ�R��8��Ä��]��-J�g+�긊��?������x�3O���A����8����U|�NLY�jc%ާ�\����K��wcy�%+$�`a��9���:���rN�	6�v\����D�m�*�8���z�kc=�R_�ӳHJ�u�����Du��s�5��E5n�\������?��D��Օ���F���=���L8`'�P�[��۰åU�(�k[�����z��d �o��WQ2�>��Z���z?��\Jb�:�>pQ��/_��?��7�+݂1p��5>�"�ح��1�ǥ-/�D/~O��^m_�)�sAп��}#��4�l��]Q���}X�oI�S��e{�}��Z93 =΀f@��#(�\�U��XaQ��f�G-b��i4�eT7)��:���/F����&Qe������6�|���x�1�C��W���/�+��a#��AK- i>��x� %�x�D5;�b�$��>�u�G��˻t�J�;��
��Z�:���e_�e�U�m�M������8A���/` ���g5�u�,�oAL>Å�w^Bj�4t��UP�ʺ?��b�6��˝�.����%���EmJ�՚���)��i�78DZӧj�P���W�)A�ASm�Cs���g�9<L
q��P�=eOk8f�򰢭�ib&�UWd�i�r���1c�-����E���˰�X��� �N�¶B,~/����kHrhpJC�*N�	&F���rx�ݩ�qU�3C����r�,=���b�s:��L�v�T�H�,�5�zK��OF�ӽ�K�08M�Ч�q��]E�F�G�׮~��|�u,��h���-�=���� )�����F)�f�E��o�^��SsM���"��!��jM�x��C��:ykC-8�z���v�F)6Y>�J��1&���\�s��a���.����o�{c⃰1�ʈ:YU�h�==�T�a�I��H
�?��%���S����/h��4���I�c�?�>E��!ٞnp���wJ~�-�ꗇ�D�.t�K!�&�{?�qֺ�9��+��u����P!my	o��U6��>��@�R����'޿M�{Z�&Zuc��XK~��C~nȒ���������^r�lGd�3�)�/6�;��`RJT6��%��3�X��f�A��X�
��c���Z�01��	r�,o���9kh���jս�_{42g~uU��A�E�gz<ݹ\D���=�Xh�paߊ���b��FI��rf�Cy����m�<݌f�w���y:/,\���|5�0y��2���Pj�����Gz���k�f����5�r�b,�W(k(��A��� �h��j@�䡣�F��z����q��^���?�#6�w�mD.�@�2�3�����ڠZ���s�6�{%���9V�?S1�x��-�h�y�?�7�B�9����O��w�IX#���
l0QC[���}����Pu�2tep�@�9�=2�LۦJW��*�7��Vյ	�}�֔
�g�f�K�ȸ�mt҂?��ȁ���=H��${�����2���M�Ń,G�Ê������=�EnV�/���ά�3%�Apŗ�W���w�qf�ֆ��w\���$)���6z�Pgd�2���}���`�h\��E��f��g��X�4E�pb�<�:�ó�f���n.��#� ���1fM�-�I����ޜO��lAi�#;��%E~�T�aj�q���POx�\��*����\-����KQ�A��.�G�f�<�p��<]"�:�����Q
�:��kZ	$'F�Ͼú=�B�Uf�A�T��XH�η����=�R����{T��_Ӌ_�#PW�᪏�DG�Q~H�'�-Q���r�:���ܵq�^<`&�ަ-�N���o{Z��vI���>j��!�
�,͸�.�7�X4�S�����h*�m:���3���&��� ����f��i�-.q֘teީH��R�S���An��kP_��78���@D.3h��kGF�ftD�����0�� :z(~��-��Q�Asc��kŔ{k.Yt�	�e��m�G���-69��@1��x���#���!���55~k��o�Dx�*O��h+b�w;�0���2��D��e�����K~Z���2���(c)��$g�
�q-09�FJ	b��mh&����$<��F����O`�R���C�p�Q��%F{�Ʒ��o�-&��u7��[�'�CPݝE�N���T~�oc�w�08�N��J��n����ʊ#��,e׾��M97��{kl}�6�<.�yڱ�@H[����[�y��qv,+�쇎$jn�Hb�3�{n_�=���eb�6��Z�T{�ĲdZΒ�Q�����%���0�&�S@�/!\���S���N5��3O�����O�<�l?W�O�h廲�GΑf�=$F�x�L�MJ�#PQᆝOCE@�����3����F���ԔtP���燇�T��m�M�_�j��3�|��t��px����^]���l�{b£-�nu�,F�鴑�Lϸ��P8�\}dTY=8B��\�]2��fU�Ԇ���Ri<���7��_ܫCC��}�HuV�(![�4�AN@3� �Z�^|/WKѠH�*�B��x�굌��}�ю1�~�Ej��4��PAT�XZMb_��P��?)Tv+Ǒ���>���T�6��v��C
/r��z�nr\��w��N�ȇ�ˎ����x�tyT�04y�o�u�8�;��J����RM�7�֡öp���I-��x�V}�~���ڏf��x��������c��R��������Ql��U�s�Nw�����:,�2Aݙ�8~n.�ҕP���n������?�F��j�;�2�S���~��噺� �`�}�}"��U� %d���&3uzAP7���crZ������i$�!BeS�Y�+Np��._��[0w���`�o9�^���%����/'�|�XC%'���a2s �t�[�����R�����=Ez(��eK��s<ZO%R8�Z�9��w�������Ì�v�}��\!K��ܳ����GC�V-�CΥf�ɞa������	 &М�w�G��<e\������~���8q��
p\�ڛ���r�[t.����8�<�l��)A,��5<_��.-]O[C��;�5�h	�z�䏫8@���B�v�D.▌r���8��'\�4��&˚G����LJ���Y$�Y`6��'|�N(ڼY�9u�V4�o�I�eW�4)�#�r�h��6^�߻����@ĺ`|��µ�A�o|0�rD�1�@��kfe�b��0Ƞ-�תwꀥ歄*�W��*�$��?�8j,�0	B�|�K���0�+�tA�����A���+MN�Ep­w�Z8�D>��$�`�*V-��B� �y� ��H��!R)��I0�W@7t*Mr[�l������/9OzۧZ �4�v���o,�����[[�oVb^�_ [j��mj�mY}�Q�y[�V1g��s[Tr�>�'�Y��p���D���&�g"�<L��6��0�#��&>-��x�Wvg{���2K,��)^�Φf�ޥx�� �W�@d��?L��/�W�żɼ��^�ᱪF�0��~=%UvG$e�)=y���`8�@2r[��=�Z�5�bo��N؇��b3�M�߹�Tj��P&Dx��7�
C����d����[!Kϝl��^�
�J�]�<o�7*S���u�FL傒b^ڞ�����e�Ug�Q6q�`�8����n�l�u�R�"_ݪ�?G�P4��(�8�g�aN�#�uP*�4��|n�/rG����#AS~�!����ܠA���� �����8���^Ş�Ɖ��sf�1�/x�y��ψ��<m��Y�#۵K�&�Q��5Z}3��M�Y���Ϸ��V�4'7���_�3j&w�	�WK�|�H�y(4�T���5S(IW<��dGc�.���UET�Ρ�cS3��^���Pq��;5w��&����e��z����AҼ��e�A���.n��Y!��������U��#��	�!&NL��upl߈�w
Vv��B�IA����g |Y��~ҍ�Aӗ7�]��m����-���$�]C�7T9�&�8y�����r���4��F��������v|~_���ߒj�����\��]�z��L��x*`&n�p^:*6���!A\������;��(�:�a�|�Q+;��)�.ٵj -e���ɉ�Ѣ�T�v��{?F�lz�6 ���u9(�'�Yn̄���0�q��)ď�O�Gi�uJ\����	��JϤ����7�8%f�/O� �]���:`�F��3�%��i�r��V�,y���Ӛץ5��=���4�ڨ=����Z��EKŬ���	�uU�w��t���5G^޿��1����\�D.���5��W��!BSɿ+���?�"��t.ӧ�����ݿ����pT+�믥�V�م��-�7�w��ҽ�k��Q�I� ���pEZ�s�OF�w�_>ぴg��0�yE|���#�hH�*�Wg���#<g~���0R4�0;\�]i��$qIz?ʛM9Gv��/Me���T֗�A�J���~�/��9��V�{��dS�,V�*�������
��{�A F|�"��sƒf�*&&[�	�N���9�x��/"�I��3��<kspLϦ&wo�B�5�@��L@<x�~I�A���Q�,�A������W�mXd��}k�@*yC��W��T�ѓ�`0�G ��~[O���҉�U��9�پ�X,x�npg,��U9U���Q���6E�u㑚�*��h�ۈLO�=�Z���D���b���x��N�����C/�z"�t�����bbs�1��xVE�3
�_�Ce=���8�)R{���C��&yV��i�u����6�t;��Y���V�dGo$�M0GO�K/$Ս+�y��`n�4q�s�d=���4�)<47��7�Q$@O��?k�b�pΰ�w���#=�?��&�~���D]BIQ6up�����K�8?]06�+��9`\ t��b�&�sy�ݲY����)��Lɝv7?P%V�P�
bu��/Y�j�>$���x��Y�\�J�/�g���6����ͫ��CF�3�.��.�������P�居A� jSa_��'�^�O-Ӊ��+�`�+b�&�,��bn`��M�3()�&�T��kr0���8:x�8�7�:������GT�K�SJ�y�t�K��.:6������)�2��N�_�_NXw{«Ďq���/�'3;['��Zt��H�j����Mg<� �0��^vg���؄���y�Ӕx�Ђ�Zҋb����|ˋ��.qѿ�C!��M����ׅ �n�Z�us�9t�Gk��8��	����w~I����>�8�w���|Tx��G\L�`��O6*��L�M#x�,��ѐ��H�e<	�	8��1�ފI�`B�lM�*�~�t���QK��� 7��[O���$�Que�%γ9R�L�`�[�m�\0^�_�����7�x����xV�d#�s�D�KFۣ/�0�F� � P���aƛb�]�/b{'�	`�(x*�3�"F�1���}-wY���s%�pb~��[��PK��I!n����eS҉j-�k5�Vh=T�kKX��?#"��W��&I1S�.�q�݌iQ�τ��aZl+uq��t����'�eb%g����J-�Q��%T,���fV����rX]J?�-��
N�6Ve#/aWo� :����F|R/�;gyN:J�q�N$�+����d���j��H�&�o[�ǥ��
�1���m]�W@Ĩh<��s^f0��Q�����Q0&v�P�y~��O]PF��^�v�X>B��Uj��=%:Dg������zC�\� QI����V$k�./s��w����0��0.�P�.��z�C�2�j��b2�@L=�ot�uH��0ˊ�e�г�^٧QV2�qE�o�_on��Y� ������/��ji�}_�tF|�I��Y��p��K�t��O�#��Ow$|3a�ː	l$AO*�>�����C�@T_7`|���M\8��;}l��k�߄�<� �D�͖��w5/�{���I4p������YG-B���L���<Y%��k�r��z"?|�e���qҍ\}��ԙUK���$�3����'���ߓ��U�|y3�2W��?'?+*.�#�X.�S�%��\sUhF���5�����1�ɚ�����d�g���:�&�"bv�Vf�Z9\WU��d,��%d�u#-]h��eLN�Cz� �a�zi���tc�%Zgj�L�P�`w�\�@��:�<��$�Z3��!�W]��N�6����6k��#����V #�3��ʕ���.�CS�:ep1�l���6���~�^����� U�����(���I�����.��;a��[�t�e2׏u��0�g�߈d���Y�XGAѝh�ٙ��)��Ad$}���ӮH6�V0-#H�=����a��Ѯ���}�hA�j_?\��k^ꔪ�?��t�6�Ih�#��u̔tJ��ݏjP#XE�g��CSh&�W]�
m��%
��S�&_66�JubU%�͔�0?�nN�9kM}/[�#�|^?ˉM�.���o,�b�P������8���{���z��O��|d `09*�ө���@R]\!�-Ud�T&!���c��Q�F�TG)b��|���-��0�6��0m���|�LB���;vh��kkW�K�u�e �Gx<��y(�f��ܺwFm��v��c<wY�gI�zT�}נּB�Q˵V��g�� B4��2�n�Lh��	��kdL�7H���f�.�a,�O�'�E�[�^9}�$���_�$uj!?*�$/��N}C��a��Z�ٳ'p[�;�r�������)у�E���aIri��py3�fp�ؠ"e�
�� �����[%G}��R����Ċ���?(�4Ш������>i\��dp°����<$����B�8^#� �����"�[��t��Z��NL9N�p`_S͏q�O
�;䇬2�Kl��6e��h���k"���ް��ù�r]����s�����;�]��~��T��j�
Zh{%�A�8����?*�A���O1�D8�i5�'I5BϨ[A-��@�}N���A^Ec�w���"Z����,�E�@��2��0!g���޶Q�Rg�7	^��xz8߱��x�*��G!G�N�^����o�qڥ��6C ��`	=����@��I8�(�S��& z�K��d6�­�ٲE'��R��~�z�o�]X�p�dsħ2��ϓn:��d�~�'.W��?|�aޑ<���R�,)Pۯw��B\Wjzj����?�m�17Ƹ��^#^��HGW�Jq�,`w������gО��MƐxq���G&�ޢA�~��jv(��0r�12��@%32��+��S3�AfHE�/�������δ��
ϒ�^'�>bI+H%��E��3LȂؑ�d`P�9��00"UX=��2��C�U��fb�A�0L�6�4e\���xs��^�t��3�����,Ȍ�����b��|Ԋ/���vx/�2�&�cIY���^�������2�ДΉ� /�!h=��d Y7�kEq���ּg"!�=�0�S��c�	�?f�E2�a�ޔ�'�{���� Az�n^�׊�u�C����LFq���F8z.�G�vl�d��*�������^���gM�I�|ҭ�a6e�迮Ss�	�Ф��*6�g�<�d^�:JNC�j.^�R�)��?���=�Da�"�7J�0xuס>��Ч��K,{���g�j�ٟ��*g�1�x�.�6���<�n�\O8��-����"�V�7^fg�v�[$QaVrK�i_Ja	!V
�Fj���x.����w�J�/4`�毉��R+��Rڌ¸v���w��[����(pĴU�ڑ��,���J��$����S$�(�1�����W�!���SH]k�W=u��o�pI!���2��	�l-���@��f��)��<����`}OW�'�~�\�OR+cMl8E��ߑ#����x�fQ����]-3��������%�f�fZ��7�9Y|2*��m�|���+^w[%@�h�t8��-��mu�;���I�RQʖ�K����oϏ n���I�+�h������9����8��[0�E�ucl��,���|���v§g��	Ӱ��Mӧ��ѩ	o��@i�X�OCeYo��߬�U��R�ᖢ���0���/��E�h��k㨭c�@7׵(�&ӧk����A OK�9�P��&���x����)��!ko�9^!l@�Q� ���+���K�.M��M=���0xj�;��jH�v�Z_�\�n9��11�˿�ǵ�_����F�|8O)������4�є�+�s6O"��`�y� �C	�,�£�C8I����V�G��^��=����Qj[�F�b�\ZP�X��4~#a8�����}�3-�+�܎��˭���/ޗ�6�oA�߾v^\�$Gi��"`~uCm��.n��(6�?@�����*�p��Q�l�j?{_���9Y �a,_3!��(tw*i��M�n#�!-˼*%�������f��J���D�ћ{�������,���I�F�YV���w�P.d�(�4c��,,�������(��sr�Lovm���8P�막���]죵��t��|H#a6����w���gE�ש�aڙ=(�����v��@��E\澼���iu�C��?s�7p2u*�GQcj��� s��X	�e 䚶��Ü��:^�<�v��������8DUD?s��2#B3 �͠[h[���S�2X�=6U��c�WQ��B}1�`�^B�SΡ�~	h��0�Q
�$$Q�����r�����TX>M�T��p�I�s髵ƞ9j>ֲ���d�K�3)&G��0W��L�o���o�Vflp�p-Ъ��/��ژ1È=��&�BDp����AV����� $N�m��
�Xw���e�*�b��㿢M0�c��%D1�ۍU�ЩH�2�\��L�+R�95�x���ϙ�TTv��Bg8�V�1=5�DQ�^�tU߹O��Qħ���s�<&o:��WO!��#�IeE	��S[XV7���̀�?�X���$)�?�P�]A��nS:O�q�\5�8���x��V�_�n�M|G��%��e|���[Gȑ|�ل�M.u�Ci$��u������Vk����cb��?T��4_D��.�*�S;8|�IH���ت���Fu��5IA�a�o�x"[L^A�@d��N���r#v��֕��>���&��r��D��d�}O-E9����E����� H���R������v��Av�n`x�u��`A�B��w]L�9�1,�-ڲsRŲ��տvR�g�_�:����*!^��\7wW&�E3v��%���t�xd��	��T2�ZxG/ �3���e; PΤز�Ok�����M��枿 
�8���d�=06"	vH?�)j�GЯ�O��b���~A*% �yvs�������&�{�����ʃ����y#�)]��*-��̂c����� kߣ�l��_��
-m�����w^�0�z��� �6���G�\U�Q:ï�Q����ǐ��K���VO���E����	�>e��K�gd�D
�O�I���}dKGVj^Ԥ�L¦l`5 ���|�[��Y؎4�I:��x�������Ѿ�$�fA�4�����ݺ�}������?�s���s�yB܉�7%m����2P�
��:ᶪM7�l�x�u.�14_�3YE�Wcfg��{�|tbK���gL�ʇ�@����s�BZ�z�w�D��3N�$�<&�`S��j�^�E�KMnhA;�!%b7e&נ����?Vg[��;�S�:�u�Gb��;Ƞ��j(�͏�
e��-��<j��O'#�ײBHj5��[�|���EH7��5�zh_U�v0Y������Q˴�ש��RE�S��$f͆��mF��^���g(OY3�=�\K7/��(�N��=�������[��p	�dM���lǄ}���Q�NØ`�D����}h�O�/ɵ~딌<��{����n����	������n�+�[���TC�.&`t���eG�h�lw���a$�h�c�%g�r�x�S�����_1L��8+WY#E��^1��'#8�t�/���oE�u���e��O5,�m�o��1����Dz\��� �Nψ9�z��q��T3x[�v�~�j�4�jp�!�Cu�����x14���)>�@{��UG�`��l�����k*�����T���=�n	�0��Fz%����V��Ϛ�a\�f$�c��(��ư��z�@�&�&`
�S�&�A�4q:�{<��le%dk���S��y, �EN0n�JO��~��������6���IU�>H���)(ѫ���Gu50���H(���P��7\����Q.8��,E�o��e���A��n^���7�b�}�1�'k�y	���u�+Ai�t���c�*�r&����� ����e�L���2�b�S�6��5�����7=(������n��:ȹ�.�d"��XO�{�C�r�)99����=J�aBӓ*��v`�]Ҽ�k�\O���#��6�_����}�fu[��?�
j��4��X�[Zx��d�+�p<e%�ǡRa3u�+�T�M�p��Ӗm�"�KW�l>�[�)��A�g���4U3S^��XM{���K41��,<�-��f3�S�=����*hD����ZF7�~�%�G�����������P��F�פ� �I-<�}���5��P�0"d�RZע����RK�C~6k���!�����j�`9S���3����d�+.�����	l	Wj,���ܴ�F�麯~�5��@��_��{�-Ɛ"n�m�`�Y�oe6Bq���/�����-��Qs���})��A��Í&"/��6Z���`w������	�0*��g&�������μ�Q�N)V�]�r��=��$N�����A��hͮ��f�&5-����0e��]Zb$��X(y"��oNE�k��t�P%����E~�S҂��j����B��,h�_��P��w�l?��9{�xN�,x�w*�Re����]�����W�*ׅ
p�tÁ�[s� �Rg\A�D�3b0OBR^�E{H�*?ܙ����P�>k��M��6�=���ǝ�G�Jp�4���rpPW��'�ч��_��GC� k�O�$Y�~�`�$�)��x6����I_� U�y6K�7 <"�-ru�R�޼8��s	�����W�Y8��Vf{2"A���0���4�K쫑�k�$A��Hx0v-��@k��)3}��މ6��E� �-�2r�M\XYbF�YRJ�_x~�6��B�5:9����{���iY��>��c'5�M��6�6�!o3j�E!�jSG[�̊t=���z�ag _�q/��`&A忚63�Sԃ0����W��s�@U��%��b�o�w��v���F9���Q<x=�9 �2F�9qx�����^����G�媊Ry��>��r1��RJ��`|��~�O�{W�t.f#k��(�T�rn}�cn��lhI�X�"�Sv�<2_��
�W�ݧ���\@B���z =��Nվ#���W��(�D{3a�\By�"!��Ȇ������H��dS9Q(����&G~*4#o@˄�\=�u��c��l��u3��(9x��2���3�����r�ݪ��Q��'��q?�o�d��⊷+��hh�pxHt���A��O�{H�V�>J�\��?���b�-L?��H5������)�+b�v�k��7s����J�4f���ϙ�u���_1ղ=p�ޙ�<�)�4��T�$�Y�d(a��Ǟ�|�yh����JP�.��d����D�B�Z�B.Q����ք��i5x�P5E�-U�"k��R�B{�x��G
���Qm���ϴ�u��Z��7�k	A�[Dg���@��/B�g^oe�|�f�v� %z/�?�~7�x����_Yf�fޢ:��J���� �Եk[�Z�ю��7�f��Ϊ�������-��X�B��M�\�F��.8=;��mhR�42�E���Ŏ���f����^�q��U�m�6;*�7���"��~9�ݹ�/ ��8N������j�>�a��)2�G��:ނ��W	������"� hz�\*�i]�4��#֑������]�jp�9����,+���a��n ?�Rݿw��K��Z��V��>��wgl�T2��4?R��ƨ�*+���@ Ԓ$����`�K�<[��|�/�����{�.9���<���C��v,� �� �,nR�է�oX��9ŽI^'�-E�yl�]ln+=t2�F�c�#W�Pw�M�j='�y���q�zNM�#�8����UnT���w_<��~`��e��� �dEx�+uF�s�h���̐,�]�{�7�c*�G��X���:��84$SC�aO��3H:/0��Z����v�ȿ&�h��aUT^��%.���[�L]�m�6�1�po˿g���S���'��j2ϯ���I �?�6
���g���5�$����{R��i�ׇΪ�5�| 4Zd
wG�aM=��N�� L�@|&I��1Z����9��u�;z�G����Dy�X�ms�R��ؽ�z#���!2t���h�������Xr��9q���-�I����n��fXa#��'����B�5��e����
K�ɦ��`eF�{� ��BA�;�Gy�n/�m�ȹP��(�FMY\��(�g$e1M(̖x��
��& a���Η�2{���D{+�U�� ��!.\o�\9>cYVN�zM���/����p��v�'���Nx�},QS��X����_ mݛ'��i���ڕ�e�$H[\Sӝ��TJ�����'_��97���ܞb�I<]�u��Mr�0�٥Q� �"�,;��a�Gq��2�"g���}��$���(`#q�|3 1m�L��*��M��w�F(�!�\�p���*�+]��.B�YC�j����P�E�:�f�3W���{�"�p�������`�܄�� ��?�IAf����/ˑTZ Jt���-���1b?Co>kv��O������/�'�o�sKH�/%y����8��	P��CrI?^Կ?���u�ݥɈ�hǚ�t`�Jr�,�N!�"���/�2qWo7�&|�w���C�������d*��"��+ݸ�"��1B!XT6˔��C��K����X���0���2>��v>ZTO��F����e�M.�F���:���(ASY2!~�{���^/!;�|��H�I��4>�0,���N�8P�>_R�=��X�>��^�@H�d\%�$o~���݂�x2M�4����E2�{m|j��h��a�{Ο��i��Q)����YI�\v�Y�o�V�����e��Ƹ���ً���E_���Q�p:>�<�N��Ls�[ﳃGUrU����M�b�qesU�q3K6>4<����! �M�J!�j�pv�QA,�`�������b�ϱ���L��'���ia�k�5��_�xx��\�h.(f�`rZ��b$P��*�6��=U^�IV�b��J���P6��L¦�2��H���L(�#�?���Χ7�߰r�����O$\��$6t�/L�77�}h����θ�*�yY��6Q�ó�&9�}��Ÿo��*95���O+)ò�SPF]�)�>V��+�_Q<���Gܙ�U��V�M���08�H6��٬�Tl8�0OD�����Q=u��^)�'��� z�\�&�q����`�7 a�TG�*s��S�;�L��!����z���1UG��P�ˋ>�h��p�v���e1b���h�<�A��WO��jP���Վ��]��`/�-�a�ECj  d�n򑏹�@\Vi��2��K �b=�)�Bܶ�i��N����#dj�h�|;|�[��X^���km���[���F틇�
�m>S TM�8#ԉ�7Pr��B�A��X���XFg"�Zj�\*��E�
��Ie����͡Xu��%��qAк��I�|Z�ܧ;�p�����D��|�83���I�{ƜVxK�8b�|�/��m�f�]��
h��)0]�Tz.&+��$���R�q]���L�O�%N�GuSاY�/\��֪%�3��)�i�0����v{��RM��8<%Ɣ;{^ǳE��l4T��}G  C�D�N�C\����x��C�4�O��nWO!��ޟ�S	���a�� ^�O)2J�G�ī�lp��� f|�4�_�6��n����o�Ck�KD�jW��A^��Ҁ>�_���AK>7?@��$�)I��Ɓ-��]Q����3E����ݸ�(3Ŗ�\����A��}�o��&�bh�sEYdN#	$y>3M��\�7��j.���|[�]1ӗįR�������Y�{�Eh/�U�oj�N��nw�8�D���W[j�yݏ�y�f�g%�B-��R��#=��j�����=��=��0��1�9!�@%�X�D�j��󟾿-o���T���w�O�Gzk�{o��,e$L<�i�:3�ӭW(컿�n��@E�;�Vx��[iS���?h�K�����y���-�x��R�,����N�o�5��n8:��$��6U��-U�>7%���/�_9�b�(�	��J)mtԫ�N#��r	Մb�fj0dĩ����|;5F}���Yg��L`Xcb9Jr��.��U�D]~5
�����G+���$��g�b!�3z�}hx����ȁ�v��
7n��j�k�wD��JK��@���P4ާ\)ru�UJ�3"��Zs	ՠy�ν�3gX�o�}Yɑ��%��"�D��z���9B�J#7Bk���ҍ
�1�J!���TLZ�{o�ɻ�u�R>�yO��6ս��[�Һs���s���crgY���\�;�lך������{��X�1��@�ϐ���E.Q�泅K��#�e�!6���W@T�E�����M
�=�ix�p�P��|=aQ ?���*>���#��͝�7`c	�ݵs���d�<T����-����'0�̂���/�p4&������Yi�&��,��|"��I�\\�?QNz*����|���6�u�׽� -_B�	yt~hj韅��;��?i)���PE��-�jAM%���vbp���C���9�Q�WS`~)�yw֮�dq���I$����E
����w��pf�J�`h�k$������qF3�z�2ʩc��t?;��=q��1��/����Ikʷ��:::tE��V�dQ�ౙX��� ��/:�(���?h��C�mmF^m���	�*�ܜc���E��N���6pq-�5�������_i�,���{�D��
P�BK>��@*5�T�F_]��m��F�G��hJ�[s���IVO�+ܷ�2ԛ�@w��UX ��ΓƓA7˓b�eg3���]��*�ƑS�N)XJ�H�*�ˤ�c,�$�P�iY�a���G��ܜ�3{;�|&�we�C˳N 70���0����6#0��Ŧt���- �$���,`����XU�r�J%�0=)ا�s�a> ���E3�-��DJ�I��fٰ��aU�-a�I�:P�7���<��\����`<�q6(��ۮ�����b>pZq���8�������N ��<u�.�����yVZ� �r��� i�s)3z����U˧|�(C)���3��R$X�����^Y4y�R!�7T�9P��|�ԍS�QW�B?@چ<���TTy��I�����x�p�X"���mr�s�pW%\Z��#��GfK�)�����xÍT$�7���Gr�ؒY6h�$�ʐO����"�F�{��`梈�Ghw����<E��O���\q�M�!�u3���Ye��p� ���.J	�S�㮳#j�Q�$xq���%I4` �.!��m3א|�b��6 ���hi��ހ�g%ġE��1ȩIsM;��$�^��`>���~�Jᬸ�CX?������I\�\�Bz���s��ǲ��ދ��֔�9DB:�B���.\��ߝ���l�$�TGF�MM5�0�P��҅���wI_���{Ɨ��ɉ���؏c��`���#��,5��`4����O���;.�/ݕ�4.Z����I�X�]Xe��Թ�]��<:�ML��A�j�j[�?BFG!s�k�Ԥ}hptV��t�Nl�C���4O`:��	P>gڣ����}�הΌ�Y�6�"]�8�"uA��?�f�`���veȰ��՞����J��p�,�:�Bx�f�1Wl	�y���)5(���t,S��N��p�4d�a&�|�D\�_J9�g��ȷxҠAn�j�.�k�&�b�f<�Q%���2�?hFr!K�tʯ��{��]TY1�Wf�>CW�V�Ɵ�^��v�3.8�i��x:�MP>�8�ǫ6j���Pf9�����`/I?;�f�6��;������Z�.��y��N��k�~`�����j:�Ϣ���M9x�5�kr;/�sUv˪ۙ��9Z��.I���4��n����J�VV��L[8<R�a`.���)����
��Yӗ*0gB=&���Lx�6ˉc�@�K�f��ꟽ��>�1�xa��$�K^yUg7�"�f��-w��fm13�x�m�r�������p���@[��5b�UG���#�*�]�����o��_��E��1#����X���G�$Pj��)��9���tr��<�G����A��|.qP���a���x�ɺ�Scq��k����3�*�V=��=�o#qVu6� >H)�;��m�ŁءW7���ȗ�(1UA���we�x�����$@=f���g�,g�G�������vN��V^8��^b�0z>4��#�2;[������2ƕ!�W��".pN����i^�KP�G��/�/\ΕD��.�,;��k�۬����hR���/�Ჸ#�J���0��LS�z�����:�;��&������������u�'V�C�[��l�Z�%4�����
.'�\�����#q\&���+��`���:��5�&R��f~mԝp�跘� �����U�ّ�|sdz��U�\�;d��僑C�y��'�g>maJr���#�J�n�̖Vs��'l֯�^�N?
�q�<����rQ�a�	?�0�
܃�r�����gd��<���l|� ��߻I�D�ڞòS��}ms��,f���Q'�/06����'� `Rd����#�C���D�'}�^*r�am������r�̐}��$��*d`�ͅ�����&�-�1�6��T������j��@.��G\s�������/½�2�]��&;���U5�G�I��[J�ر��c��V�n�۠jĸ��4��bw�,w�l�Ǫ��or�0z2#��0a�B�`ڿH��5i������������˜ٌ���� ��l�7���Һh�W�|�엮�P���1�(i�]O7-Gh�&M�^�`x<���D�ğ�]��?,��Bbo�j�l�c>) /j���:6�.Ҫ�33��k���z�(���5������W%��k}EݔT��/h؁�_,�p��ƳY�g�>���J��<���{M�;��,��C�I����Ll���;h��"� EV�ٚ��_��\ܷY|2�1�H���6cA���E��&�x��+�u*sWP�*cZ N��rV�˲GU^p��.U�`�H!5LRsW�u3YчN�C�2KZ����<�����K�(�3�6��� �揥�a���7#O�d�n�c� �D5�t�/Nf�-�:
ȹ��S󂂈��\��δY����)��;�G׍f z�mСP�-�M ����m��Dk��
�g&N!F{��~�I���!rC?wjnj��w��^���ؼDCP�#>�z��;�&-	�	u��w�MkqbvT�n�<T����~l)m%�('�	�_#�����[��= ��b�1ltD��_�\
;~�xY����U��F���佚�&�7R!gF@�Uk�J�� �<���'5δ>#�YS�
���&ܵbg��<x3���&,�.9I��z������l4���hۥ��/�vt��H�=��P�{��a�V:�������l�\��娩��cE9�4r��4�?��P�}>���҄���8�]ǥ��2���5���iI�ct�{4KR\�c&��`��v*����1�ͦPie'�����$M���uKؔBd��a�?%n��sa˴�
1�'������ rT$���kM ��_gn'�k�.G��-�����3�C�v�.[��=!�BC�yѴ�R�A�U�>̱�u�����-��cg�ɓF��e(�҇�6�t�(��b��\I��"�j���dF��V�l�9vy�!�4O2x0
�Q�Q�횗�X�P�Si��I�vs�HT0�G�tJ�A�{J����A�=%��O�;�B�9�H��b9
m��9��`�"^��"�ڢ�03��q�>��|��A\�k�;�����'+˃T�#�B���xn��������]''{��ys@���-(O��X�պ�������X��G�%����Jzh�����o��y��\�=N�d G8E����{�� �K	�6��C�ĪW��**]fDyt1h�A�)
J% ����!�#/��@�+��`�( ]��ݝ���#*r���>��LJ*��I�;�O@A�C�ۇ��h�����7������a��j8�. :����"R.��E�~�S@����w�l��,��W�i.�@ �_m�,d�C��C%Oi��@��#z�l��Z��U�8B�!��'j�]p�� |�5��#��+�����������R���"(S�TW� 51nʒ͜=�!�W��yi���6lĻ�w�T�g��O��j~�3�U{f��謃�nT�n�}�H�#�mŶTrj��V�Fn(Y$�b�R,�2P몞�~����Q�yS׻��i/4ge(�C1N�c�Y{��p�=�޿h�#lI��[9{�+`�t��=0�d(*��%���d �\}�` ���*��đ �X��b�<���n�WrG�U��e�u\{�-]�H`O>%��p^�hN!�9%�_�+���b8~�f�>h]i����np���4, �o%� ���mW�����́PF�U6i����5(����?�sts}ú��H� XÁ	�酮�;�IA �z4��xȈ��Kw�Sc@�WE��Q:I��Z�Dϐ�M?}+d8�g���l?��>PKJ+�5u��|��q�n��V��g6��A�!�t�?�~�~q�.#�\���|�ܭ����ظ��TX�I�������Ӧ��w��:ì�:�>���y���L���j�&c�y �}�^�K�ή��|F;|)$����0�vh���pBls��b)��M	�v���l��ו=W4 �4�uH*��{�]aFQ@ŋ���G)�2���7es.��yp���S�*6������x��~�g�Ȫ��ܝY�"ǯ*���D��W#aNC÷ ���u�}+����C�a�I0�@�;p�G|�2@��Ȉ�b�2MB�^k/��G�w�i�-�i�u��|F�2&޾������\ZX���x�`Fn���M�
�K�E}2�×��hF��)����AM��9;ّ̩����Ɉ9X�X���X�(w��9ƹ/��{� fф��(��JX̔X�/0o��c�2�h�������X��ȻR�e���#�������D�|�3��/P����D.F~�_�$q� O�0�Z�Ѐ���Q3aT��_?�.\������i �᜾�i�E��T��~V)����1������V[����e{}��͢�����I�4m :/*�ֲ��x��.2�4jo�g������hB��_U�Dphxd��vU����o����<-�Dmh����⭃���Odȶx��dbk�Ŏ����Jg��]O��֩�z^1.����.p� �a���V�+.�����eR<{�DC@�V��J��T��?v����LF�d��L@�+/�/���Y��L���kPe&U��]~վF�n�ɂZ���~�F~~�)��t|�E�]�@�����VŸ忛B�������E�Ā3��hN$���j�&��?b�k�贠�2B:���|pp��$W�;M��R��̣��W��*��D%��KW����}dU{�J[����A�d�Y�o���C t��f7�~������zo!Y.G�bC�v2X�/���O�(��fT\5r�ZA�ѽ�A�st+�l��`'fj��F���D���l�LPԠ�FV/؆����c��?�0�F���O��-T`�Δ�r�K*��ɥ��.�)��EP�{Q�q�>��*���Yd���s�@�6?\�B.S_�[����>X��YI^^�����{~}��G~��-[U��5���ܪ!����\�^��n�:V���d�,0�~���QXt+�FJ?�W�X�^�rg���ok=S�:�'&}�E�S���@a)&{GE�l��!�z���8�KR?�*pIT7��"Н=y���l_yp䎄����^�V5����}`�|��4%C��f�튱G]�cf�-�%dk]��u�TE��R����D�y��L��߰�5��F��'��E�!�]��rW�X�7k�v�F�ȕQ�D��������"`�)ט�{w�+"������G'�S�eZZ	;��򍋄f����JExy����Q�T���,jJm6=kB�C��I�D*0��lˌ��k{����{,I�bz�tT��L�!��U���Q;��#�z8��vyyx5���x�X/�C�Z͓�#]���W��%��q�!c�j�|�l>Z��Љ+�+t��˼&�?PJ@|����U~�3?�ک��-��@W��ьs*0�8�K����:����[s�E��G�p��&��]��H�;_�Y9WR���wx;�s|}����y��r���y�y"�H
R��ٌR��4Y�S���v�8
G$�f�~�6#2�|�?U.�ĿӔ��䍾����ƠӁ���~����C�ɸ�_�bZ�LǹO�/�]t?���RN�B�e?�(n%}�<.o5�����' ��:�Ĉ+0�ĦF�cfo�ql̈��U*Q�u3ZOC�DF�bnO]��d<�[˒���\�ۺ�6I�s�A��=ߦ�`�^(��_Pdu�t2pC�O���U���D�qphm$U#~�(H���k�Ǧ!ڀ5[w��I�;���W�i�Hts(�G[���9�*@���:���O�%{���/_4�}��TpK���z�Au����ʖ���u02�rfj,~W��u��U��3]�Z�����3(38WǷb�z��'�HM@���_!�.n}I)�;n6^k�KJA.u��H;�	vBX�b�
�,%�������$�<��V����#7$����n-���:�����Q��Â�A��v+�*OY.�1��oӱLn�\�A��H��IfywN+P�^9�ַq@�<�oXP�Hd90��h8K��P�ⵃ�ok+��U��P�@c�����L#]����^'!�r��n����q̭'�tP�:���kxqX��sS^��m�Z��Α�~��)V�/e枔���F����AV����w��U��7@t�������7�������N�a��UU�ڑ1�tgebi����"zv�d�2*W%�{��B�A}�l�ւ/��� �ݱ� b�G���Թ��W�_�(��I'fS�؀
�o�Mr1�Aw�>��v}��7��ޣ���-�Y��|���YP���7=�D^�f��7�)ꊦNu�JR��a����y9��3�v:Q���}�K��"v�?��-:S5��JQZ����d�?�+�v�����1����Lҿo�GO�R���I��5�fM����d��-��y�j�d�OJlW��Ü⒡�+��|Y������¢Q�EЇ�H���	L"�c��J /�� �GP=�K�� �3�0J�rh�q��ʖ �YE:%�$�<����j~�m,�X�)��j�'�ю=�n���S�e���������������>��,e�9�=k��<-)��M��Ѳq#R�=9 ҋ��F7u�?��[�-&e����O����S���qE�E�B�P���#��mT�yQSvۤoo��(�G��/*�C��un@:�+-,�U��g������,C�����]�ov� �D�dq��v~���!^�P�;��a�] �̪	9(���r�*�2v�A[�7A
s���K�KP�?�	����h����'��|�'kt��),���U2ry�E�7�j�y����1����}�ӫ33���~?{�-Qv��\,���oE׷�˟���ޝ��qq���K�����v��W���74���VB#��o�Ŵ$�66(�%�8�����F�x�[�D��6HfU{G��Ew6�iN�3�
��u��Q��aY�ԛG�.��t~��*���U�S��)�~��0�Fm"���+�"�i�:����H F��ڙG�kQ�9LI�u��+E#>�1�\�V#�Y4�Fg���a7^j`�X%�1�p��lͰSw#�54� Pb�CD�ۗB7s�A�9��#�5+�p�MI�)����k9�7)���vxBSoV�`�6�,s�ĩ�Al7�	;��Qs���(F��%'e�g�#Ce_![�ͅJ!��A�����L9�ʨGi�bo835�c�	���7h�w�%���F�o��%x�'�����E�T:.ɢ���+��V `
�u�9cc�i�Ԁ�'p�B�y�7�!�o�w��/
�]Ƒ���\��^x�&��)�㡳��"쮟vh�S��ت`/��݀�I��wJ3�菿?��m���3΁�i�zV��I=m���A�gf�vG�f�U6��*[��Q�U��I�,����hB�^D�;�0�^�V��z��t�;Lu�w6d���*����M����̩� \�T3�Z��Tv9�G�cd3��*�t�,�&Jd�s��?�kCD5h9Q�)�,��
e�=����E>L�Eej:ibr'�`���[��?+0"ο�� 6\<iY5�t�������#��c����6Q ^��{�A8��E]w.���ȕ<�H�E	q�������{L�t��y�U�}/�Ĺ'X�f:w�pՅ����E*Ag#^�qw�>�Y~�p_q9�,�3��Nٶ�5l5z���ԩ;z���я%�Y�fl�\��v�m��v�~���բ�3<%�J�����!&A�������-<�B@��os��\lLX�z�a�羿��m�e��OZu�0.��V�d�n���|��h�r��\]�p�B,-�ߐ�W-�4a�4��7��Ei����tSF$�x2^���0���"]�2;e!��ܮ#����p�2]�}c�����'l���#a܎ds���=U�����ӭÌII'}���ę�@�Ə�o�ـ3�*n��r=rʻH�L��~5ۍ3�뀠a�h�]��oU:�����qm ���̫�5�>��-��Dn`-�T�6D���cA�����v�b�+�
n��v�c	�a[: qTATD�r��KD��&��O/�*��������	�'n�D6
D،�����nmM�,~��$y#n��X�\!\�ԫ�F��1�<w�Q�[�TX1�35���X
�Ԋ��řv�]j_͐��S���^�g5C��!$��z3�;�7����,��5ش��,r6ݢ���$L%{�Rq)�;��H��>�2+��uh�^&M�EǄ�Uѽ����	Mœ6#߉M!$��h�6�2�s�ZW:�N��7�U�����S���g7(*̷��'8��>��F���_0
1(��){ U�|0�z�k�'�D�*~��
oFIzY��nw�u�l����3l1Q�c�/�u��Q����$��S�;��s�9���.B�@�3�6αX��l�]�B����S�V;.~8UYc�������"U�wq��R�{O��Y�];�P)�L`��k����c�a�HA\�ʥ���ӂ�	�n�YiY�(J�rE:�U],7SG�����_#*���t�����t�ny���皦0]��P���k�Ӊl �)�i�U[����0����#�w�e�/!xUȧr�	{�rM�{���i�Ś�,;a}���d����	�����c���>0�:[���G�>(�J�U�'����3gQ$��U ,�0u���7�0!�0U�{���qհa׹
E'2"p���Vv@PO���E���^��	l5!��A����J<����ۓ[44�v�EQ���?k�J��	/��0gB�)��M�_6b+5,ׁ�ѠV��:��@��d��؄���* "����M��S�i�=�� ���n
�>��8{%�6���]If#0�a�(6۞~��u�s�7˓OgHHgMxL�z�R�tJx���GSCq���5���`��6�(:l:�$x}9�.��m[�]f�I��	
8U�����+S��I�3�JՒX�,��16'e�7�O�H�&�RMM��}�π�_���R��Q�EF-��4�u˺?Z?4'��i�z@�ypʴ��.�ͱv�#� ]o�i����IA*��c�+��-�Z��'-I_�y�$R�H-�/ BI��Y?��d�=#�\�d�w��D���,�rP���j�y��
տ�%'�!�v�]��!'�g��b�HVf> :6�s�@�"g7=��]�-��*>����K�Ȅ�st�튅�A��OPLp����0s,S\��y#ɧY�$ǯ�9��X��m��g���)����8Ϙ��f���Xb)�4�I����Źz��j�	�9�73F����0j���.� ���rNͮ�Jw����h�D��S� �X��ċ����Cc�0�~�fl{ɋ�����R^��C]h=C��Ȣi�)�K�_�x(�P?pQK���EJˊ���S����k tҍ�\}�O^\h��rSA���;))i����+v7��\�"�S�e{�}`<���C[}�[�Ղh��nX� ���|����e���g���d�Ԑ�Mc�cp��	z��{v��%���ہ)6���~�0)y�Z����͸�^H����P!B������,��d�� K�19�-󂐐3[�2۟�7$6��+���㐓��
�6�0	,�U��ʨ�jd6PYd��!�X��3t��B��a3n�u�����r�	�i'{J�2+)�39݁a}�ͥ�j����]H���0�.�A�'��x�F�� �Ql4��+>@Dj�?�V���?o�����VAy���h
5�FT�6�llS���ʵ��Xʭ�77�@f�M��+7v�~� *��ˆ��m_��ºO����&�gI�:pV�J��E ����K�q"�@��Ƭ���I�,�6�g#]�/#e�CP���R�#g�2?"P/���Wx۶p���u�b�`ﶅ���z���K�J�.X��Qa�9ןt��߉�U�o���Y�1�!�n�d��|���z!���Z�b�Pt�ʕ�g]�R��~*r�BK��q������C���WL�����"T��_9�[#[��2B'��C�Q��ƿl@��|���H��X-����d�#�����jǲ�!�<�Ѹ���g?���t�hA婭ɸ��[�~/����`˟����1�9W��|]>`P�xUX݊hu��=)��?gh�!�qSJv�zJ8Gg��(Ż�	!�z����A���'7̹��Y�K3�KՇz�p�G8������fy*�,��?[L�듺�zU[+��'"�2N�j�`)``���*�s�ྉW�U�f�v�N��j�f����=p<�vGL�[��1=i��^�\/���>��S@�z^�[.n���WF��U��~8͙	�������8����#��ǧ�v�},�(�Ӑf<�%1ȸ��D��~r[��6G���o���YI4]"~7&q��dd�Gb$�dD����
 :/��dJ��G��>|jO�J�6�mG�24�Tp��� :-غ��:N�	#�x;��"�����q5|��irj�ڳ���0|??V;o�)m����CS����������1j~@��
{�)�8T�T���!b-��M�E# �����2[�Q�3%���Տ�(Kf)ݎ��z9B�y������Lx[MH�Ό�]{`�BM���1��^����FN�G>ѧ��:(�A�|�z7q��U��n�u(�Qm�C�Sr��U^J��b� l��C�}.E�!�y�
�n?i�.3�|�U��H�����[e ��)u�����
�H;�K�GA��Q��?Ϻ���_:�ᆝNE�{�C�h�s��T�B�%�"|pm%)��; ]�5��:J��X�ˮ�#��,���cT�V������Ş�t��K��U�Y�iq:���m�1��ێ0�Gfb���yPJ�[���6/��8�%����]eoa��gɤ;��H�VdB��-�ԯ�*`Q�N�	�)=�X6��4�-Vk%pV�3D|-L8�N_���|/ҡ�.*w��5����C�P��뜻i�_�=:��<�&B��Q��b	�B�4�d\���RykT~�+Y�>p�dq<2��$��= o�I�j}�G%��N62������CkNV�V�}��+Ѣ9x3,w"�f$x�q�O�����j�݇v�V��My�f4�י�';Sj����h�?�h�(O2��u_��\��]�mp�ur�dh_H���A����Oq $e��z��F0K�:-Jm	��W|��X�-�h���3��s�dj ��fZ.�r��:���7�4�}ef�`lV5ҵ�*��eS�0����袲��@+�<0�9�1#��Q�d���-b�G�KәeכnQN��v.J�##ң�cɑV�m�cI��cՂ��D� o�U�g��a*�溢����dQH���W{����G�^�<�8B.����+:z��Q{�pGW
p�F�a�F��5U�����ǉ�oy�fx�$�G�?�b����5�__=@e;�"Bu� c/����yrN~�[f����e��]\
��@��#��V�{PD!
�`�!Ć�%�IDt�=���"����M{�r	K����a��r��"WBО��{��{�yۋ�_�-<+�����u����FRƷ\��rYc��0����0�@��B/^1ͱ���	�kfn�����g�7����Ź���'=P�M�w�����0�	+�����7�ʆ� �%���G��bx-v�E gp2a6��3u���'C%i).�E�b�Hh��������:n0�C8�ZdI�g����,�"@n�\h��m᤬�Rh��Өh�爣W��NS����CP6��7OK/���VW�r�;��|�1�
e��S9$�l	㡪A#s�U�ց�&�����~�S'�[9�.��cMmi���D�� 9�%R��z�nC���>G�Y��8 �m�����3���J)�ܒ��2.�?~�F7l�U�koɺh���b�KYf�\̠�#��p��)�.�jbkJ1�f����`��b�&e���/�ͥ��5�ȤC���Hy���z��WH�_����i�]54!��[����+�R\R�-���j��0�^y��R��=;������\r��}�k�䢨 �ݒׇN��e��ʋ�N"�H�N���J��+�F�/�b�/�K�l��˛��$�b�!j2��TLj.{��:�K p�o��S6��9�D�W%��M�ժ�4R
l�P���L)�HT2
��?Ev[�4�'����Q
E�R��2�r��RL���+[
i�'/
U5'%>�;W��޽^뮛�]�l%���5C-�g�r]dʔp�qX�� 7׷�*C�M|�Ep)�~��8���k$�!!O�Ar(�5Ϙ0�wy��f��lWW��S^��Pa�JPȒ'�z���&P̈{q� ޘ��2U~�C�|v�G?`2�%v�	f�[4�(:&�t9Pǔ��8(J�	!�m)�=���N�U�5�p�!ĳ��LV��4Nf"}����a��縗�.�8 ���M"�8toǢv�xɡ��wo�����CP!�u���[��i�[=�w����c�67�r��v"�Ds?�v���]�i����L�%;O��(��HSI(
�n�N��M����!9�����U����v��d		r&.��O��_ �ڑq�ڼ<U�¢&|�V_���U�ox��c�b���mQKm���d���P��*�y2#�N�������!9+殗���j3#�D���ڸ$����w���"Q������#�t��&Eg��3����~!S��5�t��K���;�?=�(��캓�'#����*d�.���^����%�t��<����x�@1%����B��;�Tl��-���=�Z��Ѱd�)'�-�ܨI�F�CH�פ�y��K/�fy姁Y9�X"��H��ݭ%S�g���U��J�%ǀ��S�4&���yk�&`�c�	��ӡ�!�[�췂Sz�b�0m[��_!��>s���IC�]��s��y�(H>I���?,��i\ڲ�s����-��	F��?6�8�����]R�^�7�PW>MS�_u�Z1�+j�;�';�(Z��O�L���7�Q����$_�e��k�J��BC�2r��8��F��-.�����#ک��"MB�g�*dٕN�Z���.�����(1�XC�:z��F�g� ��n��|2�A��ý�����~%��y����i����Rm���I[7�o��7�O���!�K���P���\��f�1k�;�*b%[ՎCp�>VE�3��b��#E���t�5y���Y�o��ى<���1�橣�Ŭ�B�Q�)��0c{�:�����ұ82�L>O�l�S-1G�g�Z��v��G�hO�?d���(��Y��L5��˸=�ȮՓ��X�P5^�W��{�o�P�z]�;%8��M��?3�4�>��F�K�8��n�������F{X+wv{ոS� ��/EY�:f!A	GB�`ڹM@�����b�g~៌#� j����v�p41n�B߬Oȫ[\Q.�,�e�q�҃��J����I��x̓I{����npn�[�c�I�WU�l�`��D��#��R`D�ݝx [�J���Y� �!�a��>��p�ҏ���nQ-��\w&nQI��b��J#+�RQ��������`"க�7�B�!��LOϐwYem�L���Ś��5�����S�P�6���Y����V��縛1���U�j ��v�k�(3��Ef1lA��j\v�k�O�T�F��2@{r`׋���{[��PZ�hR	�$���d��K�zԒ%S�݊��jq�e��/
�5}�d����h�������S�����*x1�Yr�{�l�Tm(���1�Ɉ��F&t�h�3�i�Il$�r1\U��ԩ2�S��ǔ_�_Ƿ�N��*����B!�7�k�"ӡ���&��/l[1h@x �~�}��i�\JC�,��aJE��gu�tR�b3*[�\W�ᙪ���TʑX@��٢��΢��V��x���eK������7�Z$B��ˇö�5��ܣ$��^.�޼����e"��J�a�Ҳ�%��)|��~h=^�2~�&��r�Đ�yR����_���YY@J���0w2Ŏ"m_-O����՟H�����cѢ��W5"ܓ�{�,����E�ю!3V~�ܳQm멀O���g�~���ܚz�-��m#n����H�Ѽ��>�p-�^!w�N�楦͞.Z�S�F�/KB���֬�[�e�[�~b�:�2�5��q;#�@��;m��tcI���$-U6i���r��RB�lK�X���;J�=�8���˖�QB!�a�]���KVE�wD�	4�_jdn�JV�����ۈ߶{��y��A��+ 9��r��0�X��~�d&2}!r����U_���I��N���E���]�E���BI�Rϛ(*Ir��4�u1=��~���Bz�%x�	����N[h����YQ�D��;�?���/�ɫG�s�s$:���>�^]���F�NE�=Wd#���"ݘ�c�GjK�j�%�L����1Yz��	[V����D*TK6���TF�D�6:ևU��$���K��'���jqS��Lt�2��� �)E�);���$�ɎȬ(�v��
�t_F�G;o�i�ZtѨ�I0�o��_�v&ZBb���!VBp���
�
�4�������6zAa`j|Qxr_7M��!����6�u�(��t�9{��hp4�����t\"f����Fu�XJ�h6�fg�n�e�/#�"�Sp=�NVy�`y`�3#�)�:Ljaµ��5�����ow�-�ف�YncJn�)�Ӌ�l)� �ǟ�)���YƶFi=o�L<�Y�s�gt���R��ZO�n�N�%�Wu���c���ߨsz�+o���3j~��ߖ��vΏ�^h�$��O�_ṬQ�./5��&D-ư����8*xʉ�a&��|I$"l�A��gVc$�D�PJWŋ�֯�v�p<�Hͮbg������x
_Ѽr��?+�b+fk�(V��4_��l�5΅BI3�n$T�;��׃�H#҃�F�i��sy޵k^��E�g]}`kpEߍ�������@��]�#�X\�!�%,��x�-
�i��%��e�''"��4 ��ز�V=8��G4J��:��R�Oǜ�KN���G��8QiZ�iDܸJ-��F��{�6��,�o���&�o:y�tDd���t�Vq��zu���g�o��";0[�1@��u$�j�z4�6�~�J�3�Br��t�[#mkKD7*��V�p�j�d��*4����zC8�H�2$�9Y��m�4WGFk Y�r��I��a)�SR�S5�kM
�]و�eq~H$ǋr#(���/l���JVبV��fћ�Ac��R���)U_�1Tӓ��y=?X���<�5�iaڜ��;�ʔ�=��@�o�����ܬw�a����J���N�7��p�O!V[D��ŒD^gv-�c;G$�2c����ݱ�y:�u�گ�l���@ *J�S��;ܝWg�Ns!�t�}����H�;.e����?�xj
{���i�X����}�F�`S*>��s�%D� ��2k,[*Q�	�"C-��R���W�8o�-�E��ƍ ��<0~o��j32�il��RG���4.��Iõ����U���@���,��rʑ��Aa<�tb��፠�)�抈S�o��@Ե�\�ﺭW���V&{ر��ɯ�0�-!��{��0��Q9�{J��[>O�d&e�\~h56o��?�Y���ŸQȚ��t��tb�~�.@b���9=�p����Ҙ-�����x<�'�&=ې�� �� ��Zfީ�v�e��\t�:�q�@vj���l0DB�`HдZoxg����IG/ׯ�S���
2��<%�ɪ���75��� i��Գ������w٥tw���*�E��!�*^ʾd�W��u:���T��k�����p+62λ�S��7�0UÕ�/�j��q��z�W|I�0��96r����瓴�rui-*br�iʯ]���6�vs<����ɷS�msy����������&B]����0<����7�zCmR��!X�;x�lzt@?@�J���uGrq��uB�7�P�����/�PqlՀ��3.��,	r1�K�{?���C	Vcܦ?�~�8�Cl��v��|^��e�!̶,��5-L��Gɼ8��Y�{d�3�W�ޅ���@^��{T'٨���US��KR���59A�Sf|��1ˋ���x�+n���,΋Փ��e\1_�j�^�M
b զj�ڸ}�F/�=0q��-#�*���w����g8;�ֺ��M��_����S3��(d!���8�&�4I/p�gY3�� �PRB�~o�l���4=��A����*�+e���^�cI����[
�zi% ��Y"� �V�W��>���>��0�sG�4+'���Y0�Ũ 2i�����L�)J0�s���{׺؅k�F��J|��;Yƣ
�\���s��5R�_��gx	���W�?xm{~���	�H;�b�Qn����� HR�!ɱ������}Hv����5���2�ex�/�."�8Twfȋ�9ؓ��J�����;�3�{�	E�
��<���|p����u�F�c���_��8�4]����ǌC��O�P�t� ��G��Q�&��p��=��b$�h�N�y[n�U:�����la�Y��mS���zR�b��[�`'Z!��i��&g���[�mY�@)¸��&k����PQ7�2�x �?�!���H�������Ī��W�7�����p���sΥĮ��r�z��R��>`H}�V*.oq�e�V�$���ru(�5_Q�-"�щ��N�e�9b�G��N[d~ oH��Ldo?O��>=�,Q7�C�F��}��t#ZL��r�C���� ��&<[��'�G\z�|i���������h̡�#�
��)<CF��n���D6N*S������/h�)���^��H�#�ݴ�,�7Y
��� `z�0|n��:ؙL+
_�.��M�6���V*�؃��eq$�;�P��Z�C!�4��<���%��]s���4Q1w�����!�d��j�0R����1s��? מ�5����80�W�-�r��]�q���)O϶��W�ZČh
� ��z�+٘Ы��4��`AT�X�+�(d{���콐��l�x?���)T%��u�⹰�K�N1��@nyB���hGR/���5Ⱦ�^�3J�&��d4���Z[NkK�?������eEp>tJ�l�C�o����6��u�|�(��͹�(���������~�ѬwqI��(Lm���Q�� ��	c�ʾ G�]h�*?4�F`\��G�wϺZ��h����h�̓�4<<��қ��ɀ�r�m� ]}�@��Ա�0Tۺ�|�<��}��ռ����O�B%!#�֘Y!¨vY�;�r;>_0d1�דW�������!��%$��(�ֲ�L��y��*�b���3.����]i<Ѫ�$_�mRkz�m�l	�l9�j;�s��� ?�;\t�*��NCJ?Bfg��wS���%:�~�4t$��>�'��,�:�]���A6�^d&;��Ch�D��I%��* ;hXhj;O. ���[]�H�/t���x�q�R8���k��.+E]����W������p�d�KҚD>�uǉ��0͢�~v��YH�x�="��	z�r����$Q���r�W��}d`�9��C"1�����$(:��9�״$k� 9g��ES�z� �(�F����.M��=A�@:yj�r�KB�D�~�b�p����}f�j��������7×3�^�0wf���
Z�Eq������H/!]{Fo6%��'!�T������X%F��e�Hݔ5�z�Ui��g&��h�hy�b�xƂKVv)�?�߉����(��Xõ��U@k�@D���G��y�([��`��ʕ̑��'�.��6��=Ka|4����n��4�����������AR�.���ό�bN�%$�u՘�� ~���p&p�ȟ��<<J�'�� ʁ��ڀI����E���{�i�8��t�/�/ᱡ���21�����=d1�V+@�
�u��t�
��Б���!��+f�H��N�9�zN�����H)!	9ҋ!���2��l?-$�s뢘�D@��]�F��@M6&%3:����6V�h��W���`�e��DF�d?��}Nv�%��ڋ�Y�W��Ezx��.4��7�\����)�Ȧ�쫿��#��,5�8���R�S�PL��9� EB��;6.b�@���.L͜g{aV�&��p�1a=TB��i��B��������\��˶R}H�����H�/������޹^��vX�J�L|utg�AʲE.��}?�l&����;�l\1�hr�*�k����?<��&Ű���l��N��[��v�Bb*;ݗO���=�RM��v�F�����dQ�e_�Xm���i}佭��9@ݯ�RJ$Oi�Nc������>�Û'�Ub��k,-<e��L�*O��7�'nlL#/���Nh(�5o��2��h?�Ԇ,���t�$�C���KN1E�yz�����|�Rq#-����A���Ys�5��}�j�RU��ŵ�t��|/"<xe�IZ����T�`������Ϟ/�&�9*�p�x�6rK��b?��ؿ������?"ݬ�Ƽ��u���QF[}����w�����d
Ȋ�߱�c�w=�`�$���jc�sF���X.[�F�zpCR��$wb��O��gUR��+{*�dƸ�Ta�����i!�(1�^ԅx?	�B�a��U�y?��yv}�s�Ҩ�4v�ƭ&��]��Ǟ|�\��s�ߤ��#%w�����y�n�4#Q��)M-�M�����L�ma�r���h=�N ����>b׍�YEঢpC
p�ʣ���"i _{�Q\N�4�oևE��+��`����^��۔^+��G�*h�O�;�f3+8��9�i|��CiJ���pҏ��E�v�Ը^�������X܇�l,Q���L�����jT�pBz��ѷ.�Gl��Z�;zev7oRIQnч�S�L���e��$�2��~���T��)z�����Ⱥ3�2��8�b1u����C���T�&�G�H�5��rY1�/�B�0�[��Yi��Bq2˗��IϨ��&u�ۭ�y~̴�����@��M��G��ז-=?^ �r
!�z��nM�Hk>/�;��0c�p��#�\��7А�}`�d��V?�V�-����Ѷ�3v������RJ=!��w��6F�˟�3aȄD\o���*s4YW���c�Ĥ�)GR�Kx~HRR|�ҷ1�4#�э�"I0��]=�MxP~��L>a�$K#y������[��v0sf��ґ�]gmg3BBSMK6E�9��"N��S V�{�y���b�#�J����FJy�{�{�{	:�5NLA4���_�u��*$�BB�H��[	_�'۽���넘4"}����Y#��u�d��t����9�4�ڳ\�b����8㕿�U���H���C(I� Ú/K*��������=I1,+���Y�d(�V��K|0PC2���Ը�_s��e�H�TDB ��sܫ�5�-'!g��]m�������d
�\��v.`Z_���O��,�O�=0&�,����_�������8�Rl~�Q(R�6�o��;4��V$n�:�v8 ����1�m�B�jT�&�$p#�CH�X��V���SZf\<��b���P�Vh�r x��j�d�mםe'.H��R�����_�L^�8�nj�t�[P\f��n0����~�ר�.t�ǣ�R�c�:�f���9�4��Rjoy�*�(��},幹Ŷ�����,�2ٺp�F�D⥒"y��J��_�ۙ��V'�9Nǥ��$NyKְ��m�? �Оj�5"0�è�q��v�o�)sÆ�LX6x��o�U�����rC�˰�f>��(����j�D"�2�`�*�.2t��T;in0�P�Tw%�H�|g��8i��N�=�E�����-���fMf H3A�[<lD��D��P�������A@b���f��{:��BϧL��N��\�O痂(��E˷4�!�}�N4���J�*T�SyƁ�N�I����p���b���M?t�?�l�����;����i�}��lr<�S�������E �2�AUX���� ���T��Þ����ZWN�����o�y��s\�����/q�j�8B�e��v?@���鞯r�)�{1?zo/�W����9�F~��,��9I�uWz5#vOww�}�2v���\��2X���7�.����p��a�v��u:~�D�j ���$�L2Za-��
d� ���?� �x�p��/�mQ�r�>���gm�_!�7�A�2�琺���	r�2��6����u,03'J�p�u�Or9�����r9�'P\I�Ԛj-l��R\����()t
hU�M$lY�q,�v��:t��}`�}P����^2LG�(��#W
8'����RD��+?���g���ۡ�l�N}��͆2z�}eK�y�L���=п�;v�Q�M�c���u��͝{����I���|m�04J��C�H�1߰SM�g���<_���1�݅g�����bJ�-g�Y�Y��T^�am�}~�v��P}(,�.�B���.�L��1��� G3	c6�䎀�XGūd� 2�	[���z��3߷��u0Y���*�7�4N���i����^��A��Wk���P�\���N+~{��V����)Xl����()^��������8�aT1	��i��׬�=�X������i�%oD����aP9��-0Qq��O>~J�wA����B&-���M�}��M�2}��)�ND�ǭؓL�)��%t���"RX��ѣ)wL�3��nKy,R�Cf��2'I@�ω��c�V^��WF�9�R앴(@�%�_X+�5�7��#�����G>��Ǘo�ߗ�&cqd&W�)峕��YX�����	Xj\S՜N�9�s4��LR�u<��HJ�R�E�*&�y48D��T�(@P��Kyj�E������j0�"�xF�P��Yn�����WV���]��aM�^;�y���oyGa��:CxDl6��x	������FҸ�`�O���6@Ry	kL��ʡ�;A�0�mS�T��#g ��6�n�{�������Z&V��H���8�;Gpd@�; D03<k�AgӗY�;�%��A�mW��eN���'W����ݢ��$0b��e��=S�����3��!��V�P8؝�r��`N�h/i>�Ф����hإ���U�|��� �����	��x�W�y1�޷��P��]�K���]J�$7��a���n��vͲ��c���̈́̂v� ��j�B�EșH����1�&=�	?��G�2�������ʭY5� .f���Dx[R��f�v��腺�3`p���a� #�j��׹�io���)���J�r�4�=A8=�I����n�Q	%���w?T�&����U!5�䞕*V�X�)td�
Z��:)�`,����H�K���X�D2���n�%]�-��6�H���m�!�ߍ�۔_�U�#�}����Ya�,�D���!?�n�W�վ���ᐍ��4v���6Q�'�:����2�^Ok[_���l����1�gl���E;�Z�Oa92�^'�G^��0�q*n=�vt��/��咳��*𚕍����N�tӇBq�R1������2�<4�Hk�Qn�#�y�\]å*�YnJ�u���B�?�	&��W�"78���{�S��h��� ��u\�4׹��F�6���X� �`�Q�]x�Y)��������r,�%��2v|�ڹ�A��l�96��5��E,C�*�}�����_��vq � *2��K�D���
q����3���|XPh���Z	ׂ������F�:��G`њ3%�������`B��s��K�z�/��R��<V�X\��I����.���y�l{*b�Y鈇������uyA��B�ު��6*��خ��jo�i�O�m�9ˢ[��e�p�������]%MK����l�>ݍ��{Y�t�ar�sYT�k���#��5xq��Rƾֲ��XG�1k�[��`��h� czg:�Gȳ���Ù�� g�!>]��X���0�2��`=/����qЍ�*��F��_gՀ�$:�k�����p��;����}륯�7��<޸��\�/}��;�[�!��Z�'cE�}7�����ݱ�}��g�q��~�����,���dԒ浈��8�z�֑��f,1%WO<���y?�-F�;ʑX�6A���bX���~5x�U��x�j>�7�^�������˕�1����)��WQ���[fPZ��C􌊕�/3��+~�'uw��w�A�����U��X�Rф�`B�%'O�A�J�hfU��Zr��f�r6�z��R��r�BT�GH�Nz��Qo���惂lG	�JW�Z5�mw��F��{�+�_��e��L�*��Har~��S�x��5Կ/6 �yȚb���Ɯ���-=�����T��R�H�
��iUaW6���c��+n�MZ#ʮ䜾�b����N��R9�����Ȧ}����-6���	[=��?8��:��;�$�eNW�L�x��i��Bn�L��l�R��:<�%&��������8p�{�	�s>�K�x<��ު�c�z�5�v������	��e�,��-�N��6B��m��닟��̚v�A�2���Qd\�ͷ��o�D�c-_K82�Ԣ�_;G��Gg!�Vo�U��Pݬ/�c�|8j#=�R�ͬD0��0���ME����lT�7?�0,t�4��*;�5�F����j�7u�1���z6D��4tr��x^'�+��q􍥠`�&��,�╯0��7�.��}$K��Zy��UBY��Nn���������� s�,�pP�	Lۜf������M`͇��j?���Ol����,2꾀������#��'�d�Ι�ݴC�
�<� �;�cq0��5O/]����V�k~dA��S��_V[*�.��o���~��(�h���y��p;<�^�������|YL-������O��R�'�K�������-�!����w��-��U>������'}~)������G��1�J���|ޫ?���3.��[�nŦ����ز�B���Z�?ZA�ͪ��7��,��@��^b]�������y�2��x�+9�&}�	��/?#��N-z��]/R0<� ��V����)/�y��2�,�Rщ �Ә�`0u�^j��[r�U�*׸z/vĥ����ZG.+U5��_ޝS�5|��b�s�����zu1�ϝGAubf����5�tx�,�pO�_Y/^�>�>b��š�=��b��{oq��S.�d�^���Wށv�z�U���~Hz{o]��Q5�]�%j��~qo}�����_��(59o��*d�U���1>����g�_G~���/��껗��I�
�$���hN�z|v�˫��W����"$~T�=�Cc]\���
�~g�7������
|y�9���'j�lh�|�P��_���v��g���4�����NP��>����s�`jb
����[+V�:yN��5��.��HՑ�^��(���WW)!�w+���>�_1�Z���F�{��x�P5�����F���Pw�rA�ݣ<i� ��*,�Ğ%Cؑ��E܎� EF_
G��w��jRx���F$��%�D���TyACi������F�[GQ���H/}hu�8Sۆ�2C�?�U�;{T�S9�&���_đ=^J�:q�}]�}��Q��st��
j*�k�PL��[k	�xDƍ�h�?�:y~��&aU��sH�Y1!H��{��pJ�}x�4���;=�)ܡ`^p��F�Ubª$�#���#�D�̅f�D�g;�]E_�aʎ�&�����Lw�&o\�/�M�P��l�4٥�d}�{8�f���� �����XȖ���"x:������lGX�s��c5�'=�W�G�=��KvJ;�@�������b	�\�zj욵�`�H��c�Ԣyx&-��n�͎+�#K ]��SEd]��W������h^1qqZ'B��V��o@]�i�km"�N�+k<N;��I	7m�5��4�'�� D��# F�L�^f6�l��P�M�6k���zg��Ǐo�:
v��S!��S|�V>��N�*�Ii��B������4�w�;c������.���&n����t�>jjg*AD]�g�� �r#��1<2�������� ��ޮ��X�˓	DC����;i�&�v�Z���{x���9�e2�bc,��L#��ic�s�1�?���+פ?qߵ���ة�������U�F۷�L�
��$��d�%oA+�� !��9��V ���P�,��k��NNdV�N6��>���.@E�'�����ySp88��@��*75�ÿ����c��{�oE��d�/�9�q���F���'_�~����ʻq���#8M��5�=�a����Q_b!�U���`�����/J�>ʌ�b���}�JjD	2�)���si4
< ����g"�q��
c��������L�1 �P��Ȏ���G]۽d�����tP��N���߲���]+��$7���	��������)h|T��J�":DqKg*�Dk�i< �	m��j�E��[E�U$��b��tx��f|Y����,]���A�ϼ7��i��}�ɯ���b��c��$����ۀ�����g�'q�z��rV�7B����;��Q�®
�V�s�M0䃛����xQ���_� eӰ"�DJ�/�J�A�ooL�fk}�E,�L�����џgK(��0�s���?�����9�6i��_�_��4����$Χ���Da^s���EV��<#T</�>�V��P�ȡDOywYSS>o��]
�x��"t����_��%^���7�6f͛A9K�36ޢ7�)U��� pu�M�NE�8�ρ�Μ�ည^W8Ǯ	��k\��g_w��E�<�Râ"�(alnK	zCT�{��	<���!9�@���E�f峹�*T�Y��4 �;���>ݿM�Q�H�E+_�n��P���Ң1.��<{LFF�,���&`M�.��I�p9cN0�&��t������=�6';����g�e�����=޻*��=���O��^fXf���!0�J�l�"�%�k=���������fj��p �'cX!��3s�Gd��8��?.��fW�f���$�cr���x��@%��c'��bH~5��b���(l:�W�3��tE&��.��y��4J�l:�j��mi�QG[�3���^��c؄q�B1+�Hhx������?zڕw��{������ĝ�x?P��}�M��!��Ađ@��GH�z_I�/kGh�5�T��$Q��20]0�-���n_�J��7Y+���ÝQ?�HK٪1Y`��+��J�IAM�nI0��;�mR�D��{G�����z��ə��+H��TS�	q�[B��7&,I<�ϧ���<��OU��_3�'���ag�0�c�`��pYqɕ�	�0�*�Y���:� ���6?3�oW�'�{��u5��b�\��,�Ȟ�`LBM6�ugm�7����O�R[)��i�ee�S'���ؼ���;1N28r ���a����Ӓ�8<r)�Lm'�3oPq��j�D�]GO�A�y~b�|�Z��~�@���#�=Xy33�*T^ZL���i�UQ�
��$�HF	��Fm� +�A��Y�c�#�w����F^����6�o',����N��%W
:/
�K���%� �܍�a�����A{7�3+|
f��q�Q"W~K��5�)13��e���q�3�N�1��Z�iQF{�33#B��a��s�	��la�/J=�
�|BDW9���R��c�{s�"�*У�6�ʱ�~S�'��3_��)�9}�G�"��m���DR�̀X?��8r�J�!ne��$�[WS��,�+b)z
��6� ��X���l�6���5;@�^�\.B�D�/���&I~����N(j_^�6���ލ�CTp��a�Q�Sߤ[�E"rG3�\.h�l�k�G��!"�Ɗ1�P�n.b�с�j>�����};K�"猚>�@�����b]��Y�HԫD|'B{�`0 &�Gι��֫��kL��\30%B�N��+�(�=1�u����ۼ.��A_a�4��$��3:m����\����?���~uEn�B�E3i-�)'��'�m�!��թ�{��8ĥ�SS�ݳ4lZ����79T��}TH�T!�G�$7�L!�tߩl4h����J�d���8��m���Djx��/$�خ��C�b�*���4�é�	^ɿ�O����4Y��n�@Zg��8��m����J[@�4Iڪ� B���?��~/++0Ù���4���/S�����
؂h܌V��?�'�k��t�⋴���êӄ�T�(��-�J�Aj�6���:T��ܶs��st[Z%Ծ���ǁ�p���<	��]�]�'x�ljp�s�����	U�+��d*�v�Y[���iheɋ�@�#�@��]�S��®EPԼ�W�BZ�j����z��x�R�A_v�C�*�\�g�~�dH-� #T�q�+������O���F	����H�������B�Z���T>���!����V�p�GnM(�#�#XM2 qj8�f�w���yu�jC��:�nw�]����b@����6��ꐮ��Ct�=��ML�{��FvE�ق��>"���H t��;-�q۱Bizhu�[z`,&u,� %�X1w�RJ^+/��=������YT�'c�B�W�du�L��nj�չ�L
�#h�_EZYg��k<@�$l�;�&���rD]�G1h�#����%{��%YH��U�W$#�w�f��D`�-.�c�O\��ӡ>���byA�S�p��>ت�!�R�K.Л��Il�E��u���n/ՏoB�chL�4�h��s$���ֹ��"��﵍�S�>:��E}�lf(f�3��E�0�GmЯ��K����P�����D��G��l����d���Ci����m�r�c�H뚅sf�9�H��6��V�4|��;�,c��;�鯉�=���_�r�YdW�0<�y�>�Ww�H-�wF�cx�X����j֢��&;��ch�$�;�}G��m�2�4�푧�*��x�.Ց�5<��H�2��������L���w�(U����Y!�����v�ClqcBD*��P2�͇!l�J�u��{`���פ��>������*�y�|(����n]]���6�`��REZ
;��8j�����@��$(��	F\�Ĩ��.���f��N4����Ψ�B/���΍�PA�"y�-�Pv�?�-����@��T��3M���;ch#�4�O��kd��+��a�=>��7-'"�_�NR����@#ƭ�y�_�%+�df)HC�q��.��J�)������N�"nWƫ���f �B{��_�|EH�&�J�%TKE-����+H�OR��vB��?�cE���;�)�sㅿ1�z�14����%��*Qw;&V������u�%�=Zy�%�o��ͯ=�����L�����#�2I9=��`� �	�Q�"蘾� �<��*v�Or�E�:�m����a�<���+�D�[��������bX�I���������O(�tD9ߍ^�~|��P%�#u��"v5�b��藺���2��\�)nF4�:�B�	�� h#����%��K�v�Xʦ��*�X֞c�ZX�
��;�6��M~�Օ71FtR	�].�k���v�&�B��\u��N��P�`N���MI�XBN0O�9ay�,��2qM�@M��߭jx�?蛷�����A��<�ZAL�3���v����`{��S7Ũ(�#P�̒�'�LT�Bn�9n�;7����݆H�N7��t8w�5�� A�>��J��Q�b��g'���3���S�X�p� ��,1*u��W��g��7K/h�.�P��)����-]q�(=El:0�Oo�C��K����7������K����B��3m��F���4wؖ�� �V��!�ͣ�>c�)Z��%�Q`~i�56I)��w�+�0k3��9�
��Q���t�l��N�pR5�Qäj�lyS�;썿�8]a�C��4�<5��,�G"��7S�
~$�\�5���}[���)�5~t�p�����_�V�3�^�~��:��o��B�VY��.���3j>B���7�$@␴K��uw#�9[{�>���h��a
�"7�۽�mn'(�B�Y��9�}j��b	r!*b���P�,E�v�P�BɈ耳���)�������"M-��<"����r����@�Ie(z�2�NP�*o���=>�D.�W�����"F�E;�.�����5��[/Wa	Ȏe�����x����p�Q���Mx%���S'�o(�_�KV���MpY����ɹ<5}*T�E[ZJf.z��'y	a�l� D�>Cʒ�?r�6�GZ��h��2�F�������~;�fj▦�F6��OL~��d$�M��F�J��H�c�+�¦1��#qڛ��'Z��������؊uI^�*q�ܑ��ͳ��7U���O�	�N�6t0����"#�=EJ�7'|�5�<�~(�����i�{�}��vc�[�B�_��mbL�4\\���[�e>�5h?<��� F<�V�T��3��8���?-��!|�F5W���c��uH[΀���T�W5��P��Iɔ�����a^e�I��m�C��<��_�h������1�*N&��_9��;� W5��il��hR㊧�f>=��`�]1Q���P���X�Aٛ�*��c�\]J���~�I-�R3Ǟc�}��r�V��%��h&�?\��1>�ڔO�#���t����] E/�V�1��b���*��������%t~~ڢW
��!��|t�[�5�Y��t.����πDě���>��|����ܥ�@����>�3�B�q��4{�j��t�1��RF��^d+[#9������-,����h��֘��
�]����؆zPku�
j��_�Z��̋�&�d�8�mCd'[��=�4�8���g^e[/w�	a5{�ug��y`/���\j����`bo:ꪑ&�C��K+�g�-�rU��/Y�����N���;u�6���Stǥ/
�S�K���2��P��SH?9�$C�0:�\����m_d�ϣ5j��kAn`��_�Y��/����ړw�<)�Xzޚ�n}�(��b�a\�[ڸS���u����>E�_Rɿ�= 
3B�%)M��X��+��xۘ�1��꠵����9WH�_�օ�.�S��0���f�G���}����i�#���:�bGq�B��T��?���!X4|� 'v��J�Z�=����|m�@;v���U���h����6�]�����˿"��o�c�����ٰ<B�2<u��h�:��U!�]*��]���Ep���j	�M��#�2�D@܊=��^����QJG6gĴ�/��&)��4�T�,a?n9��C�r��.�.˴B[6������yˁ�\���W�:���E=�l&j�t�إb�����A2��z��azW���n�կ�#�&�t�58��P���f?��Aa8�CT���Ċ�����u�P.�b���tODW$�X����	��m�Բ�n��=�Ȇ���vNDB�'���x��7�W�n���4*�e
�;�~<���j��ܥρ`���$�����Z���od�?�+:I4;'ϯð�/p]���vY����_����X�K'9��M,�'�jwL^ȃ+�P��@Ko�x��a�"[ ��f�jW���g��|oI�F�(�a	��\�?��̶����z���R��{\"�%Eqv" (�|-r.���$ ��'���wo~����I��s���<4�!��ׅ"kd�x<�U79ѩ�w��̶q{�Z��Qſ�eV�d��r?+ʚ�2#.��H����2�uU��ObR��6�Fۥ7S|�{�#7�܀C��?Ҫ�D�cO��H�,:��E���\Xv�s'��ݝ�e��d��-�����R
F�?��{�n�>��;����<��=ΰ����Ov<E]���]�e��S��*�_�;�czfܶD4 ) �à C��k�3Az�.A�As7�����|��6�Ӛ���j�Q����I����LPeԟ�A�AT���#�ωX�ժe��~P(M���{�/
����!.IZĭ6�-�?���#�\�^"R�#�m���>J
��ֶdQ8��w������#�~Ǯѻ�BPg|B.�QƢ��%�8>���BC���Y|����z�j�큄$�<8<�)ԙ���ˌq�?Q��TLX7�aF���W�]��FpX@x��V��]�"�Gh�����Iɐ�<Ѐ��Q���?��O�����E����?�K��,1����T�9��S�|��M�p)�3��#���!ł�
,j�@_�c#l�Ўx�!j�8"1�j�&��1/!����p�Ƒ�&v��Z*�ć�}�e���G�ܡ.R���P����Ģ��'Z���0��?����Lu��,�d��ʖ��Q��^�!}Ӿ�uKd8S������R���o"߹�U�A��m�A��5�#5���W�U��� $��}F0}�`t��Hݴt��A~^��P�9��������6j�B|r��L`qR��hƚ�9-�ǯ(J�G���
	�?\�ˇ����`!������P��þ�9�XJx���b�	\�
�Υ�=�k_�' ��S��<��*ů�&���82��?�/�){��\-�'B>��%��ڼ�T͉y^qʷ�`�8`��L#X�K��9� �/�D>�p�� �He�SdZX�Z��F�