��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�����uK~YSokj�&�9ȼ�P������şd�rU�gb�nEg��e��`�"9H�bLr?\�JK�߾�Y��WU����4�UNvz�URec�:�Ծx�B;e��烡�	�a	�a�H"����,��Ο�z���۩Xc� o�ѽ�F�IgRb�A�~��t_\�v�b	 ���5��G��r>��T�CF�/�ݸ#Ɍ�td�M�\FxT$��٘��ߔ�M�"�䮤�Mt����  ��{�������]������
�P8��z��c���b�S?�*K��O�~b�*����}��f^鎸ݯ���֜�%�	HڧX�Pe�dҥ�1(�2�S�Z�o����}2�<�w����[�j#�>���wNn{@D|ߒ���a3�U����g�;'G����t�䨥�x�7��S�W��sw @a�G�*>6�t����5�7=���6�_/�3�%��1�:vZ-�^�)G杮��:���m�&Q��$�r�QN�!Y���DYCz  �GCd�=�Kb v�/ ��K��&P�7�:��P���$���.M
C\�jp֣����B��(%`�x�V�6�ߘ�hvF��ˈu�QhiY����ȷ�w�n ���U���S�q�!BK��^�8v���������ۍ�X68\K��Yhb�pA��z����bj�$���(�� r�3�	dy�"`��
䳨A���nu��M���GК&qG���~����Փ�=�V��:�>a�T-���-�7���pІ�95ֵ��m0�6��JKԱ=\iӌ�X�k���>���K8������,&f�_�Z�Y}�r�N�Jlo,K�W���ª0�t�z!�����λ���xJ�I*�����ȿl���D,T���ۈ�l!�'�#��I�~�t5Q��pK-]���ttB+����lS,w�w	�2��oW<��@7���`������Ɓ��E�n�50<ͽ	��Q=��K�:N��4�v�5�I�V��%��N������hM���F�����d�۽	�
�����*������rh�y]���g�k�&��񾕤W�q���۹G�1��#G���z&�d���i�N��ъ���v������/�8Nڞ1|w��yW1lm���鑗��D���q��^�l�U�*zf'�Jg�WI�HX#k	��mi� �:�9`�%����݇�a�t55]M��i��a㄁���XP{;�_��tb���_���Z(�����G����:$�`�H�W����c%�=%�Ֆ����?VZSz�j찆�������qCBI5?_�m.2�lV+d�1�J/x�#�J��-k.��|G]�:t�"�t��ە]@>��%3#�����b<�:�I�X�Ǥhr�I����sI�
�O��HkV[4�G��>��z)��v�������(���'c������� t'�{cd�����`��@�hg��5d��:��=��ӳ:8{�g��_Q�1��&N}��ӆ'F	�8(�Z��p��7u-|��J����m��8�s�(7���;?��� �2\��&z0�2x���L�@�0oƇ��=F�66�x2��UV�~>֬�^>GHAD:��c�7�ּ��5�-h�4x"��k�2C�E����b1����Y�K���
�㔪Б�m6ZNj�3��0a����L�Uf-�l�~�N����N@ s�ȝ��d'�I�����J��1��ı���u�~��ᕇ��l��Eb���x1��J |�rf���&�)�Dx�T�`mo��v�j�=jD���,�h�ʰ � Q�5�9g�#�z�k�#1M�������R�B�m� G�7�ʙ��ؖ����j�񵵉{{q�ZA�`χ�ړ ��p�w#��还�-�rԭ����h�۷AG~KS�5���	c���u'e�-��z�D󋐤� ��#��.S	�9"a����Ǝ�䷏YE��Y��n7�i��:"�n�P�W��d�(k�d�$=ʙ���Pj�֍�{���پ�f�����>�O��¤�r���,�->��ϸĔ1�u�P�)򴀢Ӡ�O����ۿ�����B����c+\��D��T6�>-��8�xXuX6YA�R��v[¢=<[��$Vû��|0�ܱI�<��)����^��/���q^�
��@ĤWT��T�G����W���;Ӏ��0�ֳ�&��ҹ\D��|��X{rn�5P�n�O��\����B��8��1������!և1�3�'��^}����"a|�p��������@}X�[���=���-+\��~8/S��r�)h� s�<u [�>̴V��6���6$o�G�y r�Q̅�g�L�Hڴ.�l�2��C�`�u������+��M�lòlyP'̝����A�!A*��I�nC���A�y奇R1�7a�-�z�-��
�;O	���-s��A0	�+z&�6M�ZU��`)��Él1���_��룠��|�<!�v�޹}�u��㨂����]�9c30�����sn�D6=č�Z�Z� YE����v�"^�b1=jǹ���V�Z�r5����mu�N'����5|G�<9R��P׻#��5��L���~�#��gi����ޮ������`�C�����0|�|��m6nD3���R`����0���+��0�)1[�~El�&����i&����@K�`LzM*)��c�}H�zm�3HΩc���U�j�����V�4���-���6���6{�^i��[��	�� L��Xr�x����0�h
�l_�ն9�?��1]3ĸ#��uٶ�odD<��p-Ё�����l�m\M��%�I�Jٮfn�x�R8J�qQU/�g�/q��x&
j�;�pCcd�af��fz����PS�H
��SZ~�Gy��o�v��h~]��*������}�����|���gp��x:u�j�Sc�$8QB@65OB�]��Uy��e�t��t���$f�T�²�����,��y{x����8ښZ�V�����Lu���azb�hfh�2�C�s��gWɣ���Z�1I��3e����)���5|�]'<!�v����	�󯯿����(̈́����P��j%�۴����mb�a����0w��s���^�E��e_5P�α�6��0_Z�5���-�ܚ!����s���/N����ҳ�?�=,k�AF R���h	��b��+\`}�`Y�\cky'$��?� �KR"�w%��OKHH��65�U����*����[��\�o�8�&V�'4vo��V�Uob����0��
�l�N�ȋ��wưp2yQza��"�q?�
O0u�2�Y}'�9i���B�^v��1{��Zk_�WsE�ٯ���X4Y�r�>b�y�&dm7D��͂�J����~&Q'��gǍ������B�^���?�U�K�'��v.�����E'�r&� ���R��Wn���i)LR��MB4����F�al:�����it#���a�!i>?_�8�ًG�����)p�Pgt���N�;Jh��ᜃF�N*$�lA�F&N�G�%mؚw��ϓ�8�h����[A[Mz�Y�=�*"���}�ASoUd��W";4p�Da�t+]f��Z��-k}����O���@�}��Q�"W�' aAA����R��#�Jq��a,Ռ�z�ꖻ_�������>��������r~��_�C}u$0�zro*a�Ӄ.=�M]}\��}~�K�<��eW�5���/�̓����ݹ;�h&|B��9V~�]�~�#2������o�dJ/�LРs|�/0���ў��[F�/�	���{'[aW�?"�f��k1>� ��k��U�q��P� �j%w����b��U��Ǔ�I�#��ENq��o��f�ؤŨ�+Z���z�f�W�攳T��~+��i�qYk�v'�)C�}o�0�	���}��/=@��&�ٞ�6�����'�/1�A���L�/�F���b�P㐵��O��7�{��oNxG#����v!�W�j�
���T(��,�1�1�;�	�p�D�4���h�k�z�GG}�ێ����Sh�3�1@i
:+Km��-b,t�yj�O�&��ǲʺ�+�<�:��:~�5�PE�.=0bL�d�Z��*/���{�Q4.���V��8ݝ���]XGȻ�>����rʵ��it�~��o��V��	C�jW~��0d�f�Z�����Yx�~��π��=�
T�o��Ƨ��3�~�����?T,�;d�w3G��y�~3��ǘ�[��+^���!W:P�3��!X����[,l��~����YT�W���sJhUB<#�B�h �wuM��L-�eɫ^V�P�$~$!ی���ʈg��i���*	��Q]�Z�z�KK|�H���c�{�j�v���ǧ��0��"g)��&:5�3��ʗ���܀�׈�q�S��%4�����<˸2͐r��-�$M�ɻ�Q��2���r��	`w1,,�8\��7Te�Ɏ�$Ⱥ}��fJlN�[�`���m\�r��T��x�Z��5��?�o!��=<Ӓ���~�z��6����ڥu���8nR�2M�~�k�Q��²F���;wX��S�GIyk��*ð�u��T?�5�d��Qi���7?�<#Z�V�s��i��K��^b��+����]xrwS m��[�0s��_�������?)�����J�e/`����!H��*�f�2gq���R_��q����ŵ-k�h8�I�ڄ�/.8a��)4Ro��B)38�΢�4�z�w�!K{�L���wC/��mt��a{o*�ܽF#������5���f���  gΔ,wH�������f�Q��:S�<\z������}�P,��C�*�m@A����D�u��bl��#�s�/��/NI��'O�p��83l��x���nP����6d�`MR6��X�_�w���kn���N?rt�=i��c\)x�(�>��v�Z�$���a��r$��C�s�bM1�V��]��6]<扂�ѝ:0�m�}�뾺���n{,��� ����]1`�4�	���5�#�߯,m%@,=���la���Y����_+����Km�9�k�,��6�0����sB���+o̠�!K�M.��1�1���a�޿��Mw��'9�O[�����{�!(�
B���A@+p�f&�T-N 2$��Mw!г\�]�-�~����e�p{��kx@�W:��5�|���W�A�Xn�2�(P1u"�!g\���܋c&��/���/��[:�x����^mp� ˙��4�ꗉ�c'd��Ʈ�7��>Q��A$� �����r�^�� ��;v�"g����};����`Ԕ������ؾ{�Y$;-gt[�G��I$ܭM��"-��r�,}͟�ob���E�����G-�=H������!pt��5��P�S����k��N*{QM��7��K�n�W���#�S\���%�Q�E5�[H�D���9ū��ސHސ�BlRD�"ZUXV�
ls���|��>o_�[2=E�xd��N9���DB�|��2nE+zV�%Å��n������;6�����{���<w�	�~u2���a$	���_�n+�^5,�����+����9h��A�?����ĺ�Rִl�� ������qZk�m�����~%''tkټ[��xȰJ`?�]\Ͷ$huyؖ!��65�c�=9�Z��r�(]����O.%oF����6#�� #�t��)�g��F��Q����秸�J�4�F�G���ڑ��@���bUq8�
t�	6�u����[i�WG&a����PTG��ce�1�$O�C,�6ܔdg@�e�1�?i�X̀��o�w)+-P���02�B2�n��[��6rfN|"%��{`�愁A���=��&��,B����H�o_K��uO���ˤY�jR��(m\���"5�؊ġ��RX2������j��Q3��{�,�	"��l0�v0j|W6׹�i��ga�2#�"k����pΠ֬#(�X:��)�hH��=�L[�qo�I0U�z��5�X-+�_;;٪�]��i�����N��Y�=�Z�m���z`��3�bl^g���$ �Q)�1����M�%@��O f�3[�����C���Zk�$Lmn0�������3c�3Q=��a���"�B�O�F<�v�`�]�U!��U���8�J�O`�<�G�D��xd��Ն��M��/;ú�cG5W�n��FlO赦��n���6��c�Q�)<3ʘ���2�ʡ���i�;!$��ͽ������ʕ���LiOzGI��M���g����g�j]Г�Ч9T�Y�2�'X�����~ h��D����P�t���c�����2���V�Bcc�g>(n����eL�M�'1v)����}���Q�*�g�R.M;��02��5	Qy��ƯB�~���	��Wst������3Bm��	���v�T��b;�p����D�v���z\Ұ3���aϦ�CK�p ���|wu�ϑ>�]�빮"�~�P��~2�r�Ƨ��r�6�;��M�Po�6��̹�:�{a/`��90��\��b��VII ?��t�@b)�W�� T�p�}e��Xa��[P�v}D~�!�������)�@dy+�j�}�D[	�-��(��E
��=���8���?�����)�D�T\O�#��oxw����Y�X������Q�K�y�ŬAܐ�,�5���{i������F,}���ō'�����2�}�c���6�80r?U�y�:s�J�7{8�-gPJg7��a��S�f�jLy��&���~��ls`�l��
_�r�QΘ���'�6=��
S�i@�T�n��S��"�$do��'��`
[+���H�`WZ��m��FaQ`���Z�<M9� &�$�'RW�H�w�s�Y�3c�Y��}����0o��FR��E�/8�Ry���9{��6z�Ъ���:bA� C� _h	q ��|�ӊ{�����ޫ�~�voI�M-��7���F�*������-���`{g�4����X ����OU��4nh�Z��ןBS+O�_0\]e��Z�w�˅�k�}��hc�t7�|��©��Υ�"����1�z"!&Da(/����6c]�Ł�V�TӷX�9ߦ�C�\kv4�d��%����m,��s��Z\���AN�WҺq8�RQ��0��G*�#�"�F�Q�a�2��7�j}]M��9�����X��O���a�1Pܠ�m��4�9g�`�#Č}�����Z*+�]I%��jT@q�gm(Z�!|�W23�T}��$<�S�K��c��ѿ�T&J�_9.g A�%a�zx���X�^(-
B��}r��)8Ÿ�qfL-�k:R�>G�~�rC�#�������G��=E���p��y�8��S�۲��{M�Љ@F]Qe�7��b�����ȷ��ŵ3_R�����v#`�w�_�h���T�4)� ���X�+�E-ëJ�ɐ��;��"�W�T�F��P;��'��'�F��3��F�9h��i)F�N���VM�-Mu�Z�`6,q�An ��u$2������r�Ğ�I���T$� a5����� �Ɲ��qAX@m��\;�0���%����i�ӭ�6��}�(���O@�G,8A�ܡ��B&5�G��b�`}\,�o�'�Sf�:��+�������ڃk��
k;���Q�1)��FD�V���᱾�t5��٤�/N#�iyR����f�O]�Ӯ!�O�?x��?��򤉹q��2�����i����^%�9����4�!ٍe;�����O����:0�������\r�Y�)f��k35x��?�y�`E}ˢ����➟����,K��l�ڭ��Z�:}�o�)cC���/����^s��ի5e�y8_$�F5V�����c��m��^��	fCF`�J��l�ΘWh��Ri������b+ኖ@{�DꟘ�Ҁ~��-A\��*j�S��$l��g�E �;?�������T��E�-�P�T�U�U��#[+������0#Xq$�Iz�v���W�C��QH��eWk�b����U�
�Y"啵d,��q��ţ�ӱ���l�T?�S��eK<�0d��e^��-��&6��+b�KP�a���w~Uj��L/�{��B7|h��Շ���'�1�;ʞK�קC�����0�?�Nᕨh�I�����&O��j����זØ�ʴ;~�����&T{���T���Q	����<�b_�	�i��9�����w-������#��z���O��@�=�=S	lv�i�5�U�r�39�_���ي= ��]a�U��O�[JII?�
���������RX�N�x�� F��ṕ�m�X�+~����y=S�Udwֽ��1�_0�m�P?�8��Rfz];��U^��~����0����Lz�u��@��l�/-�;��0���,)f�)5��v��d|�����}��O]\Y�O� &�����4ʈ�1	͆Bn�/�V��?��^)�X �o)h1����@R�?�wh��#�j����5��H	FU캡|�˄xt�Ρi���#E�dw`��a��I���ph%�A�x���@$���p�H���b���+�,}�G�
����fK�}�7�.r��ݹs�K�So�L	Pp�)��g�]C�g���y&�y+G��L�tL�Xkʢ���@ E�J#�u�0,z��;�iNe�����Ih�; �ǰ��#��a��g�W�α��N�_�Tv���&QTu���ݒ��pQ�Tf�ʆ�Q0�I�sκ�@M��n���
Iǲ���/>x(8P3��`�9���^��̒�0�9K��F�ܲŭ|sKk�N��NY��~��J�MBow�Tr�̩��ʮW:L�w⣩��)R�'fy#�HfVWb�gb��`��T��3�"�.d��/k�3=�$�X�<1[�
C0j�E	C��	}=�{N�?h� )C�ѫd�͓�gC쳽�Z�P���騅�g���x�������Ќs�I���`��2��)w-�L)A瞪�d ����)`��� ���"�:Y�M���S���}�7$���xAq	�~'4�n,��>���#%�����l�뗲�$e�K�|��4��2���]��<��{���m�YA��<��9Vr��$Т9n!$b�R���ȉ��@�����A$��x^5��)�=�����~nFK���葔3dY1o���$����^N�̫��`��5�0�@`�O͐r�~�]�c速���ܡ�X���<<��X퇖?�rM�X�Th�4������V���f˳o���g�W2{{c|Qy���nq��x,n%��F�@o.dA?V8=�*���~��z݊-yt���m��#۱��h�"� ���L2y2S�L�L@tnB5�i��q��� v��̯�s���u������S��)S�j�C�"zb��V�G\yC[�Ƥ{�tK�UD�ě�8�
"�vCy�t����z��;�w;J��G�/���ut��(��x���դ��
�m>��54�*?q���Q��'u�]��@y�@�����/S͚�i��|���v,Ν{ӣ��w�Sm��Ɏ"�p���.��H��ݯ�7~����ٟ7ϙ�-�҇���ͱ53 #!U
�8|�呍 �E��ԯ�ł2\r�ڍws8�F��
.�&�=N���;3���as����p��"��W�� rg�e"M@��YC��1�w����<���v�k�#g!� [�a,��2J�6���6�7��&p�ƣA��[r�MRi����Q�=R�Əq]�J��Q��r�5�*2����U;�őc���N���P\���6�c�����H�ŕSb0�?���Tkk:��:1��Hoo�_|�U�GZ� ����U�+����\M��+��Mk�fȰ�xA��L������1��fA��'�JP¡P�L;P<�f�̶B��
�gr�\||��<0�~����H;r�������9��3��v�� ��M�g�2���w!� 8
�ZN�.�i���	whAWS�7�l┙i]B��D���U���(PĎ݄U{��ӏ�i��>"�GߒX�d��H����4�9��Y	+��Ӆ0��u�&dD��Jz��>��w�QN�4S���;C��S��sD�O��L�[qaN[�CЎ@��v��ؽ,��s�=;����v��Nץ�n�`�j�(�,�L8�����˥%켑QHU3�l�L�X# \N�Q@,ZG�c;=S���հR�ڿ�ZHΫ��45�U�1�u),^[N�}E�7�!%^K<�4�׫����{U*�#���J�@I�a���/�����:�hc�p�sR�ؗ�
ӑ���k�l�/f��B1��ߑ�{��%\����/V�6�%4��<�e�~��]��S��{=l;�e��M4��9ܹs�~_r�3��~�`���TS~��Y����Y�B��xc�g�ZaK�+����J����jv�qĶ�-L��įSK�X����,/흍� ��s������;����0$PM{���gYf^���Ȓ5�id!�_1���xJ��`�������Q�� �'�u��r䲄OQ���"kZd��M���)�f'�1O��#�Ld|B@dia|Oq�O���g�lGt`��E :�Â����>�@!ꁡ�=N���CY�?�%�|)�����a�S���o���k�.B�֩�Fl+�)�<��g��=dO�M����Vjn=q%���%�NW�V�.����H��ۗ������m�^5��n�_����c�$�$�	LwO�N[�%c��|���qπ���Pyc���N�u�;|jK�A�;z�K�P��[r��7������}@�XS��a����e7<��	�Ձd69�aX��V��39y�9u7����SV
zF���L2a����䳹6O��c�&j�ѕ���;�'Cn�V:X$Y}���D�4�:NN���ُf�@��L�R[�o�{�� [3��e~�k�U-�������xp}4��"s.�|x>):#���4E�I��_���X@K!G#��;�W�	�w/}��!R��D#��EG��h5� ��
�oMZ�a]Eg{�sjnh����5?<2�H�˨ؒ�=.��2]��e�@�q˟!X�����_A�UP���,�XsY���"�DG����=3Qu�wЁ>��H�%��̘���Iu´�·�/��e�]�d.U_UvW,�ƹo��zY^w?�V������(�ǳ ���h#&�4*����Y|�c�i�>�k�k��^y<I]AE���ǡȾ�C3�*�7��z0Vl'���T�_�T����������6%�F���=�.U��@�����2���sʩ�������hZsg.�>�t�K�'X&G�[L݄8�YɭR�Ak���_��&f���
��VKOݷ���F����;�ݘ��h����6-�%y�E&��K��K��Kˮ�j�H@�fO=�J�T �x�	�x�h�����c�
ǔ��W.?�|��~�������V(T��"��(�.nX݌v\���a��Mڡn��
e��9]�q�:b✬Nu�h�[�^H�pLVpi+`X.����`�'��S���3&��u	1]z�b?�}%�u�� ��ʼ\7�t@M(���6��J����`�C4_�դ�=��V �Ci���t�x7������������ys�ː]����X�jB�%�/f{x˦�V���ڱ[�(]��i,�T�ά�ɥ�2	�9,M.���p@ S����S�$s-��B��4�r�����o���Pg�.��V&�\���v��`����-�.��hB�9������_�V1�_3���ȕ���r第f#�V�f���nB��<i��l�t�1<Rb�����'�=�Ǭ>ry:DF.;����a8�.�1�P$5������Ѐbײ���s�k�CM�t���V8p���2ot�:+�{�FTLO��/wIc6���Q$Ǣ��@x����?�V�gm�5��pŅ�.7�i��塣-�B�V`jz3ϼ�RE�Z߂��f����҉�5�:!{U��<��eg-��B��58���P�֪1�'#��XI�$�r�}F��i�槀qF2-p��o��.U\g��>�7��(B6��,��Hf4Ј��c��t��U[�@� ������!�<R����Y�r��:��e?F��}l���uѦ����ꏋ�a�Q�>�S�^l��;D��1w�8���,���Jwt�H��
����������V� ��	��4ٴ(iH�7CRp��j����e ��.�B�b�p�#��!�O(0n�����`���W(�F�RM�d�
:����RУ7�J�'ˉ�����8��l�f��=O���\f�&�%PzO�qB�a|s��t�	$�]M|�1�ն�2\{���|i ��6/$r��&�<1�7��8�\��9������L��[_�
%��ƶ���d�hGD�Ҥ�&9F�k�:�^�s�B�PW{D�v/h\we����%�ⷱ�94��W.���B��S:j�K���M��~1��~.=��i����pJ7����� ���M��޵K�%���՟�+s�c���h�j+����:Rr�دL��A�i���;����Z5x���,L�|3Y{�ѿf�e�m��M�<���$$�[<�}p�+�U��T��T��Tң��(���|�8�a�kd���b1�>��7��";6#�0�7�p[��Sg�߾�ȐG8���@���% ]	�,b�����V�S1���SJ,v/
�Zx�Gxl�q�:\کX�@+ƪ޺5���%mR�t��̺�p<�ID<����rF�d��j�����%�u��>��#�?��Ntɐ�}�m2>۾}~�M���:Z��t9i&B�Q����W��dl)��Y�����C=��b^)ئӉ6ZPx-�&7.�UV>[�$�9S�WF�)hJ��s�'���3�¡�sc_��e(kX9Ȅ��'�i�J�"];��(�V|�CYWn�Y����>HN�.&�{3��tĖ�
�x���֩Ƶ�؍�t�F�	��	?[l�Фޠ�"(q�Ϛ�D��J�[��ao�A�f4��Q��ᩅ߄�h�
v�#����d�,�R>)����� q��h��3��,g?V�Ht�α$�_�~�9L+R�i. ?Vӯd3V�GY��\m�q؎B�J�f�W���eP.������y��+�
{��g�q������g�
��8=�Ճ8�)u�D��F��鳾S����7��f΍�jՕA�⃙T����>��!8��H���w��X�l�~I���[a`�V/�k���~R�J�[���gN��]CS�[E2�=f��S�W��Z����W{����6�meq,�uT�Ϧ�����g�L�r���l����r����_p�`�J>�n�s/�A�;z�Z��TLY0h�����h��z>�t�S��e���%A^����j�dȽ3���UW�@x���� ���]P#�Ҧh�s�ޤBܑ�l	i�9�sCN�B���v�8�_{�W�S�/t�\�7�;ڊWY��ᶽ�>����S<O|&��V�t2�5y�>��Q���+�"1�X�u�ÝA����cV.�ȫ1hbf����<����Oͣ�ת*�5]
-�I E,���� il��k��������2a^�(�w������|7��������n������brN$_��WX������gc.* �f
�-rp1���$@_�yb�z�"�v�%�m�@�c0�<���eR"�E�0���}�`m�&�/��{�(�I���W	<�i%O>'ӎ��R�� ��%�ѫd�b>�K�TWo`uh�&���m��ȸR�,�Gx5�l�0/"*��Y��B_���C�n��k�x;�LY����y!����ѐ~Q��&��A��V������O�P3	�ro�US�͖�V �3�`�ځDeaM�������Z|���0�!��i|+^v��C���z�{۫�y�ꬥ�3SW:
/"+�i����������/_7'�3������r�R�v���9q,z�}�/#�#��q
��e;�j���Y�^� ��GG���E����Q��D�as���<Q���Ɛ���yp��� �E����t��he0N{��qq׈���@W�+K����ܭ�G�S�̿2�-� ��3��&�کQ�:��)r�c�Y�z� ;I7�9��@Æ6O'�Ø������b+P��4#�>�#NH~1F��Ȃt����ʕR�n�[c���ƅ�%���xyI�S�ց�
LQy�O���F�V	!7��v�\��lM��I��=:�K�ڟ�����a˥�f�c�B�p�*��L��U�����G��2��BG}iR�Aj����FW;������+򪇊��ֿ'<*�؃�D�v�<���lFݷ$���zr}�8 Ii5�x278lA"���%Q�u�sf��7� �������&�6և��Q����"�[��VnI�T�A!��Բl�g��-�T���n��Zu�rm[�����y;��1���h�^BK&��T��ݯ�H�Ku>Y�WI�4�� A���n��n�z���v� ,
�#���ϊӅ�4w~�}��k[K�{U�I�َ$ �j�����\ ef����$5C>��I֎\��9	21�uY���X%i�lN��{�e3�b�1ߔVvk�e�5�u"���-�}t«�ؙC<FJ�!>4-d0���B*�K'��k^:��C��[k�ۘƙ��6���9	�}��Ky�u&�bl.���Ke�T����m�}�;�\ ��f���=ub� 浀����*�(���\s�	%�3�=Me�x�*]�B�탈A��0�..�|�������>d�$���!��]}�)h�Lˎ�*V����'�*;&9���mA��jVB/w�:��L��F�ދ�ɍ���S2�*��L���\� Z7k��_���q�O�������7�����_4�e����(��L?��k�;P0��'�w;O�\�/mF��������U ��H�����O��UOʞJx̄��j��*vp��8q�5M�F���1�,w҂�tV��G6:e��b�	{�lPd ��k��W�=���Ɠ�Sp�˞��X0P��7�'9�~�A�wp-�3,��&����z��O�^�.��ݮ=�`T
��c��
�u���B=�i�M�P�vSR��P�C#b�]�WS�U>�2�f��Yޘ�:�ə*ęx��r���!c^���=�]ads*�a������&�`���e��Oҿ�J��t�>Is0kV�uQŒ]��N�F)J��I��i`ⲹC���n�'�wC*��d�Rv�f�D�JE��4Ayl��ʼ���X����q1T'C��Y2���g��c������{Me��)[%�M@s��E@���n���U'ć/ɰ3����7����zp('��1t]��_�:��^t��Ss�2�HSm���vs$���p.�!�M���o��Z7��e��z2��f��A5�e���/�[��@���;�K�u�kG!��f<���N�w\�5>��>��m��j�E�}�/�`�sǠ��]~'o��'T��:}��V�`/f���C�^*h,au;���tA��vjJ�s�D����S�$uV�{�M�pkvZ����#�=���A�(�)����7��>��ͼDǻ�I���B��v��c�q��I�|"�(��֝~bN�l l���4,I z���lB��V����+$���U�\�!P����������a��Z������t�������o�X/h�����4�#���Ӊ{��f��g�DQ
c("��5Ou6�X���坅�.��].��j�����Ƌ>+E�iZx2�0_P��Y]���iU�׉\kS�:��X/�]��9�k��#��	A-n_Fq҅�Ef���<�@�B�|gB(�����(Y��1��s佃'���/��PB���邟G����ʰ7��#u�\M��A�..퓭�?k�]c��.�ۅ_������N�����^���B�Tq�|Ifs���ld�����P�?[�Ð
�bj�B�A����C|�<PLw�b&5��ԓ;�^�r�w�Y���y�qk=����0ݫ���AY����xb�61�Y�\2^�-SK�NN���U�x|RO#�PQ����)y�л�{S��#��$~�A;���bT6�	���VO5>��	�2|�|:e��=�>eV)�$Rw;����=��������w������}�����
7�2�|���h��߿�DV���7}�ޝgW���]�+���y��ˇyɇ(E��X���iko
D���Ė����O:��-P��S$*x�i���[��C��Бl�JEe��'����}%�V�6�S���]Ѻ�����f/�#��'Sq$?���z*�q_��UGRҼ��m�� |T�b��[I��%:F��L $I��pݴ~���>oǙ��]��M�V���MkF=���W:�������:��Ϊ�m�띅�H�t-�ni��Ki��`/��^�c�g��>�j��T]�� 3�n�h^�W�j�8Wd�:�쇟}�M#6���78౵����*	3Qӓ孏�i�gg���J��)��]����Q~ѥ�)j>~5H�PJ$�˥O�EZ�L`�Ç@�x\D�{=�D�c?!Z��s�S>aJjq�-A�_�	��� �&�=�����ve���7�~���YqZ��*�Y�|��q��G�6���DRٙ�&��D7�2��TҾ	�S�d?ie����j�ȣ�� r,���D �S�䂾�*���^:�i���A�%�##!���N�P�qh�x3Qk�xۅ��X�Cw�Ec�Ɵd�r�T-�jO��ް �7�5�&׍��l�P�.�MA��/�L(J�Ɲ.k����\����P�|^��z�"�!��J��
��M!���V&��H1�E_P��(�4��j���I�W�y�v̋٦��0����g��,xQ����1����%<��흎���]�1n�5�r���-:2��]j��[|a�-Nti��R���3����͵:
��H��" W�G�si���D�_N�d��׭b��n{���n�.Rx�[&X�����H��1���+��J�{M�3��U���V!�v�.h�c�i>H��ٯy�s��Z0@�9�#�OV�N/c.��Π��j�>\YXϠ"�aW�ʒE���EgT��WCq'qb44Q�$"�r{@ǔH%�-sQ�z�Eoi�J������)Ws\�7���b���N+)\TP��^�bɯ�δh���k���o m��/��$�d��RX��O�_��#��%�<�!�BT=$�V�H�4��YW��Rgv��UOY󼢃�u����;��y�b^�6�'���T)v�Ǣ4Zǹ	���)$T��I~C���a��0���ڰ~
�n�T��У�*S�c iՎ��tܤ(e��O�p����ςd�M#i�*�G��5Z>It�&�
�<&�egAE�8+��fG��wʊF\�*Z��q���/r���-z��*6e��L!5\�WF=�U�P���(��}��������~ ��l�"p<F��5G&{uQ���UT/ b����C��-�F�爏�Zr�][t�^�%SK(S�=��Ȏ_ɣ�/�Qm�_���AJ���@E@'y�u��PM���$߇r^�cZFV�(����"�悡\g-ӽ��Gd��ud:���b�0�/�~��2�?h�Eގ\��p���/�U>��%5���V��](�al܊��UD�+(ӄ��4��UOX�Ar�]7l'/M-�J�J��i۴�@��^A�3��*�d
f�y��4:�����H&a���t�� �բ!%3E�����)�(�e:J�Zl����;�vo�crA^K�$B�4#����G���찃P�!g({Q��ńG�@ϣ�p�?o�e+�\��C���\:��Ka�Y&������j��C��k������g䍼�X���?� D�X�@oWv��e�������h����I�b�GD���WcJ[⟤�b��\4����e�����-'d��"���m�)�L} \W�e���h��!-w!�6/R���,pH~Z�͓��1܀��59 �p=�0z�AJ4m(\�T��So�9�ijQ�!ٗأ���\��*kof��T�z�n��E������/�>�9O�r*��>�[$�X%��Dw�M���me-�l얤��h�,=�A�'�Om3Y�ߖ�B�#u��)�K3a�I�����YƵs��/ -��"�Z�A�;�e�M-\B��T>�%��2smBAZ×-�mHS.A��8�N�?Ή*��"�����dcl���;���j�����q�#��5��F5�/m��������J���4uc�������0�C�PtLv��֒Բ'�4���_L�%�:��?�����O�A�����"9�Pi���V���S����/�_MMU{#(��<�A:�w�/���L�hV��v��=�O�K;U�����u���q�������٭��VU&F��5��2G��J'��T!�z��1jϙp-6�@[BY-�`НX_*f�7צ�:U~��+�!���2�Cq�������(c����S�6,;�r�d��,����FSN�+�I�(�93�$��>gU\L�]W�UaK�䊟�+�o�͘=7��U
��iȐJ��
}~�����k�ۀ���]͕����P��L̽����b�@~]���cZ4>���
��nq�/&0�`/���3������H⥲T#NE8�������6
6�������,�)��pR	�k���!@��3���)��|��)����Q�(��}\�����#�e�e����a����Dk�\��^m��Om�$[�:O� �\��vs�V�髭�KX��S� �ʪ�ΐ��c����]Lb�}ꢿ��h��@ZZ�C`b�֢�ؽ�%D�uW��sʾZu��U�
�j�۳��P����(x�Ʈچ$�~�2����\E{��kZ��9�����nl=/0����,����r��}�В[�C+a����L���d�U��c��ѦR��'����V���;�����I,B�wH�C�%ר ����XS�,���E�����0O}�`�!�/�z�H�n�rz(Ǧn2�t�|���KsQAK�����
~�Eמf��`���6��n��L���K�2�X�H��)�I���ã�w2E7�s�2���t�I?�%�����<���dAs� ��8c��b|�������D��pի:"�6{1�K
QH�SZ�.�����S����X ���w�iF&^�tR�D5����ͯ*��*�s��uj,}z��M�䔝�L�Q�ņd�������*s�R��a?�#d�	�f�)����Cv\Ǥ1��+h��}�=��'�蝉�'���ٷap���MG�\F�����<�D�+/>���j���
?�� i������DB<VȈ�iM��;�XP}e�B�ѷ�ya�R|���@�mM��(Jј7���yU[f�q�ol��dIR���JU����nV�ν���"�X�b����v����{�V��%)>m�ȿ��*g�Ng� =��q�h�ܕ�Dm��red_(ToW3Z��UF-�b5�| e>�`����-a�1䥿Vb��܎�����2�����}�-�������9�<ڎZ3ў�j.-�y�$ejH������a@u'}�^Ï#�$]�@5����B�~ܽ]v1�c�"���Hp��*
�/4�Q�A�w��8\]�^Em��
Ϟ)����6i�f��ň�m�($������b`���
e�9�-q ���q�Rs�<P��馌#Ϩ�Вf��60IO��̩2L�;�I'�4�[ԭ���N�L�"׸|��DA��L��z�v�GV�]�آ����1.%�iD��IT�s�\$�"�t�����7�(��]7K��F�{�����ĥ&��=�f邦����.���^����d%-���e�j���Ć,����N�l�u��L�*i�:����*��>�m�% `'й ��KZ�,�D��-��gM�B�\U�Ӈ>����㤀wE��#��s~ %d|����:��9vS�����#����=�s��1M�A�������0�ƪ��{��?D`�w��w/J�b���M���}W��o�Wg��&.�l1t�����������y����왃��������� [���P�I �VH�%h3o��v�E���E��{1�:�)]ji<6����{,�8��i*�4;j��`k��=�`���;�i�B��p��u�S����Bn�A]�ǾEp���7\7��Z�x��?̎S�ZB,,v(�y��D���� {L����s>�Ŗ�Y��^?v2+��4ixg����*?R�߭JTG��
�Ǐ�Q�\���>J���?���8�#']����͗
�dIf['�^珔N`��HROv}�+z�� �,�y����h��L}�]WLіGr�M]S_�$�Č
�i4-y�p+�ѱT�(�)XG�O>��m���Me��*l��A
Wp����K(!��r�7w6^@�w����/��U1W�^bw���:Uיg?d����ˆ�GG3�����K�'��`�^��7�R��1y�x2\�Y��64��J�9&�qa6��Q�1^O��F�ҟg��̿��ĕ]nN�,mn����*S��;s0S(�M��˫�8��!��( `�j��B�_wÌ�j�}�v*4yGMb�E�ϩ�Z����ޮF��cB1�58@a���g��*P�?��a�:#?�0O)�7��N�ձ����#��������.�Q���6-O�ARoo�û����b*�Q��D�r?�y�],����.h��1�;l5�1�U��YBb*��\Sڢ����1�S�?*�!��|5�,�xv&d0�/��rx(��舥64������y���Y��M:���˂{a�h<�G��c�I��Hhxj1�	�����j�kE?�_����T�@�a��\=���:a#�*`Zߚ���J�t�0��������Czv7�%�o�7� �t�6�}V4�x��n{k�ǌY���S[vQ}T��o'�=?{�$G�aeM	�"/!N%U���i7�`�|&���m�>��[�=�����Q[I#7��8C{��a�u1!,3#%�4e�%} �T�I��)�L}�ql\n�P6b��1�6��D�f�VS����kmaQ��c$�b�G�,�.�\�
��&���o���=���C�1*s�&#dq����|���<��n������z�+mO�S�R$ˢ�F8��l�m���:�< �S�WWΘ���
��zeF����74�}��oG��O��~Q�D���z�0�	w����p�F&nq ����]�=:�S���SwS�f��Q�dK���A$A�u:3��)��Z�Au�@�"p��s���#��UA�n�&��a֊�`}��P�U�4�Z��H��B[�D1���'���%\"�T�O����*�*�Q.	��l�$�w!�F�S�\A&� {��c�=�;��0g�\#�&��<���Pϴ;��V�F�#`D�И�d�RH^V�p�L�e�������j*��G��o�d,Y�ȡ��J�'��d�UV��p�����UZߵ�O�׵��^��=�90�l��gc����ɍ��5�`�Rv)��Xm�4�4�RZ�����O?�O�t�<,�I�ߊ:8��m���R��LX����B��d�H=�v$���s�4#�ӵ�W)nKR��Q�I� s���	1��U��&0�c�@�M�q�=�Z�*@q|f��^�
'j~���l%w�{AI����(ȃ�vG��'$�s� t~)�] �Oz/��V���ob�^A���lh`ϒ,`��������1�1%���2�4������킭8�δ���I{n�����;=kJPɧ	��%(�Ҥ-�1�h�N�}�4R@4�I��kr���^�ޗ���B/'�2Ԏ#�@�g@ZgH��J�X��f���8��F'5F������Z�Mys��g>I=?ȋ��/�6R���ݤ"���ܑ	�������]�$\@�c�S��?�BYc�N+
M�(��Lt���/xIݘ���I<��J�����!�"8\� �P2ȉ���C���D��=��4�Aq����%�r��y���Ca�fλ�2���7@��x �!;�w��'������q����\��:4kD�R����/X�{8y�ʂ���7Ԗ�u����&w��|���]LǑ���Qh`�ץ���M{��qx@;�#�Jh���q����6�ܰ|-S�ز��q,�D��y:g��^�˳�d�0�]�xd�3�R�O Ff�R6��w��S�Gw��I����崺�x���Df�6�������6{y��Hkg�uZ�4)q ҩ�q�;Gj�r~���Ӣ��ȅ���pА���7i�C���A�N��nl���q�	n/�H2]sP��[�������+7(�3ɗ�`+�����"�݌n�D^E{�̷E�qU*�1?����7��,Q�|Rp�֔�͙��h8�8mNݥNi�h�)_]��`qqf��������,���\X�\�
p����3.x��NO�-^����N���Ƀ��gƂĆ+tn։�F��@�g\�����v*U���ԅ��ILK&0-ΨA���(9��$'������{Y��d�Pqo��m-��:���t�b4��{mw�jR�+��!� ��LЌ=�~�����g�����kͨX�߁���d8�f�����p9�W޴���b�d$���1�j������'�u��˓ب�^�]\L�$`z�`dF�sZ%�ۉ�OG �D�)�C
p�\8#(OeOOO�s^2d�:��è���l.O��ؖ�0]�<f�r�T�G��(�����g?�eGĀ��D+�fMε���8�ypXD��G ۀ?�;�f�ӂ�~e���2���tj!#�ۋ#d��zc^T��ǹ�:?��$H{�w`ih��Tyn�GL{Bh2ѻYM�֒����"FݬN��EB�ub��`+OS����4m�I���/�χ�rH�F�0��6�^����AF�J:�ɚ����L������l\w{a@U�m�1��GB?4�S���Á	�/,��D�7�[ݮY��:6�v�1b\RR@:_u����(�YFk��r��%=
�&�Q�	9t'�/"F��/�U"12�<(��UQB�5�������P{���%Yt�K�Z���Un���d401m����z��ma��e�3���c�	�z7)�I:vQ��u�� ڻ'F�Tݳ��.Z��%d��su��H�O��Ȅ���۾�W��n��"��\�����)���}9x��t��0�:���$�A�B���B���å���㴯�\ v��}�v�5�ꉜs!�٭ ,E�~�4W���"��.KULo��fK��u�l;��U�P�#��`n�y>ͯ�ݥ��+�M�������[�f83~��/,vn�+��?R���3-����n�#
z����2�0���P�ZW�X��4�	g~�j7�Q�Q�n$�9v���Ԧ_߭b����Y.���;'V��]�g��B�%�kR��D�qqG�F�R�;���^��:��`y����U3L���n���t1�/2����0O�^_����n����~l����	��k(u��y%� �T�9�qy�(t��K��n�>����~�dl$�c.�4g��2�,�p`(�ΨZ!MJ)Ցҡ,ȣj=�XnN�s/��d��-��f�G)w�e9?t!�D�9��X�lIL�=�1���{�SV����aťL�|P�����6�7ծ̫��� �8�UA�ԅ�TO� 8����B�Xw�f�(ec�}m;�H�?��U��Dv�����Zf�����ݺ{�F��A�5\S���Q��e�y8a�� 4���Tt�X]be�l�c�l-�oL~�t��OM6D���k>��l�V�sG��?y�11f��X=A��P��j�l�迖��ф�af�\q�I��֍D�p�d|�i��1�����2��_��N��������`�C�GI0�bPc�p�N��*���|�/�q�X���"91�ڣR�~3���Ո{����mL"��V��-��d�*�K�5�c2�XZC��޸�B5`�����/Ny������=p���� ve�	h�xX���WL�T���Y>I3+�0w˚��j}������|���f�� ��:�GA�$J�@��E��c���_>'J�2+���)��[�,^xsJ�ֳ�,�mL�i w�/r�~�����$o~�N���zQ��JW�AF�p H��A�y��$'�I���a�%&�za�H�}�/���8t��3�'� n?�1��˜rӰ`w}��	�,�	��=T���-c�q�0��7�Rjx;\�%��;��?d�{�Mܟ{���Â��wU�ӧA`h�S�\�!o��/>����:�h�7(�uI��Z �
A�"�LQt��6�N� ��2�x�������Bq��#��"yU����_J�A�J߽���3�U;�i�?��bS����x�g�_��Rp�<�?�{O���f�|$�?�:@��)Fx7��h��Е�	P��%jewaE'c�Z��I�E�>�A>�}=�A��f}�*�q��eC�5��%bW{��E���~���d`/���)K��̿�?�=�ܚɳ����[![��c>ϑԾ^�|b�4P����L�ǫ7B+a�����2k�*�7�>ٓ3k�]Ƀ��-�"ED�r+Ұ��uNy߾���� �6%X$�O������_���<������Z� iv!	��/&s�u4�A�$��7�c�q_�1AT9�$�k���̳@�,d�Ta(%ok�w��)^$�����p�I!��Ծ��Pq����c�f��M2I>0W���)�D�G�>��𞇑A�"�X�ڪ��ș�Pe$hШU&�@M6���rd�����#XioN�������i%
��j.Sst��G��I������;���V��#���;�%��h��?�j����l��}���+��eD1��������ly:(�W
o���~��� �r�$C:��nQ�~F��ߜ�'P����4��OI����=�k�FQ(!5 ��θ�Ȍ�p�g�žh���DPaHR�+��~�W[�Sjh����	ђ��kZ�@-�I�3�v04�4"��lE��ps�x��)w�0 �����"��9^E�{ǯ+������Ӷ}W�1�o_W5%{�G6U��t��n�	�.���*��~�uy<�`�)�+�����߭�*G��ht�Z��O��2ao�^��+>6~�s4��͕j� `6;.e�>�`�He���� YDf!�0�}[_��G/Aw��[2�'#�&\�_� x��*��Hˢ��4�P#Rݾ�����
H1ÐN&���M)�X/՝>lt�z�t���
fn2 ��Ѭ#�����Ì���������T�T����8k�Hj�;�1��p�8���*���'O��ٝ���0�z۟ ��Z~LɅ@@���-\υ�Υܞwo7�$�$Q%���́��
�%G�g���P�U8!Ck��ٖ?s8
�{��$�t�md���7D�V���0�g/T.���0`7��Z���$F�����y�7�*�	l�ЙӚ�}Ȥ;I<<����6{��)2+(->��6� &>Iv>��5uNo��U����x�A)Z闄0q�hq���,��,�ҁL#���Ⓥ!3��K	/!�o�fiC8s9n,F<`CIϦ��z�rQ�ղ�r�z��5��w�kYO���,��,�i#i@������Q�T(�j���"N��xh�TQ�ȟ�hu�$�#��â�u����/U��8M)���(X���=�7⬵��$�����Kb&���;�����t�*",q�#^���L"l!��-��zуEO#�Fk)�ɾ��6Y,p�]i���
U��Ml��j�h��?��l�1i(>�B�ס�՚	fF/��E��u��j��|C��J��9��K�F�b��03��c�|�R�L<�+�ʓe��{q���Y�$��ߩ�>��hn�Qjȗ?�� N����x�T��9�;92���i��%�6QP�/\u_q�+��Se�p��˭��<pxH�)��v�H�5�S*�����k'Ӟ�d� [���;gM�+y��bw��鳄	O�����== x���2���%��?���ſW���i$��p/�G9Iޤ�e����p�o���Ѹ�N0}�m�Wq��Q15�ps��lSr h���?�e�`��=���%a-�P�r��D�iH�����8���}�9�Nuiο��~�����sfV:M����S���N2/(7�;v=���cn'��d�.��U,�5��H���z�aZ�l��������Ē�,P�?�7�J˥{QI�����/���-C��[�w�GYhX�Oض;�q8
G����ڻ��+�f�]-O�������w����K�G����/J�T���G�>�)�ό���x��Y�AY��l�?R>Ȼ� d.Ӿ4�T�G�?>,��BT�;�u׃,ن������s����{���}w>�(5�(�͏�9���П��y��V�Xv�	dY!R��z������N���aJB1����t'��@�gv����VUg庑O����ڼ�V���w~��A�.���2��lկ; �T6 ����;:qYW\Ä����=����y����&�P:��k�)�y�Q��$��g�p*l�������`T7��3kΔ����ż��lx:\	�[��Hh�DO�.Q١K�l��S�~��J.C�1�,)m4�6^�t�M ʳ�SNJ�w^K��dS9X�'*S	i~���7 �z+$��T���z�T�����<(��a̡+��>��>��8�9y��F'f+�t���!��T�dɽ�Hۄ�65�
?���t��a,��`ЋVIj;\�B���R��h�N�\��e>qR�jU��v��y>G��E¦��DP��w���k�'l���'���((xQ4*��C$�6	���c���nv��q$���-��6YrJ���s�z���m4.����vд;��4/���*�ύ)$݂�E���h�;���	Ü�1���`������1\�4��ڧaX(�[�R�A��!�<�k��0a�\&��x�A>w�j���$��˝�ʘe��c{d�4����i�������"��JKneIv��(1Q=-��%���j�Ƌ#�󸂹�-�r��qr�
"��I9�VJ��@M�Óƫ�t>,�F��v@Xz����_���Q�Y\A�$��C��?��Pd�B�y�h傲�4��
��rs�sh��Z��a1w�2�6�K��ʺy-�ŭ����s�ާ���A��A*��UIP��Eg��$l��b��P@'�Wb�r�O��rV	��2���sR��NI��t)"�Ќ.�TGn��?��W�27�4M�)�����+�#z���k��Yr��&6�y�f�2�����9y$���Vz�F�gG����c��9�qӆ� ����69�����Z�M��f^��&3�����.��:�c.M��� 7�(�mM	�Oj�:Rױ�RscYA:Ƅ���ˣ�,�ޯt�y�u�'t�:Ma��>��aX�r��0���9"1�E�+��h���Yw��y��iX�|�ae�PX�U��u6|2�2��#Zl�_�1�J/+�DMt6vBxRCj��I������3{��Ą��Uyb�}!,x�<Rє�z��u~�ֻ�c4e��m�D�!�ż"������3�Õ��4��\gw�'�f�b+��A��n��7��'�a�S2�b!��2!GU���d� EYk��E���i�r4��b;@b��v���;�@<�n���Ê&��@�*��kX6��_,�	�l)�
a�Ę�#�$1�Bg݅���3���ʡi7k8�ɉ�^I=M����d����5"�y~�)��{jjsU�F����_�j�<1ݝlz���*�ў��"ĕt������U�wrv��7D��t�.�o������� r��+�#�t�ކ|��3���x+��/�y���B��m%��M���l�@�|�9w.\���0����o��.�@����0"�]r���UH�����?��W�/��/vV|��6~	�-�:0^�2����~�x�3'/�GkdD��'Q�Z�ɐ>�c�l@�ҭ;+a�>d��y@nT��u �g��,ԥ���x��yF7.)�'�o��o�u���~���G��.ʏ�h��d����`�Zis�{��i���0�[k�?�z��ɜ��,�-�@�M��l�I0��r� 7�n׀$����t��7Q�Jy��F��	Y$䶝�n�1=?rآ�ʈ�Ȓkԩ�����$�m���d5�1-?���W���a�-�\.	 �\ʋ�0t���+�B���U��m�� ,s��^���CkTI�G�ڸ܏����  �0ڥ���7��Z�"`�`�%`Q�����Q��W��/)�P+)v��Z���?���~@�}���,�1-7J����j.�����[\K�"�[@����%�nk�$,C�;�0�������
�:]����dU��&�
�ٟ�"z#���*���� x@ׯ�(��af�۪�
j���Rw4r�I��Vhh��g�����0�'\|�/�NɈ�X:i�(�����f�=��ں��$ҜucB��Y`p��z�6Ag��{��?aS�R�{�j�����EH���a�E/%�V����0peӶ�햟�� ���%{qB��J��*Oz-?q5a�dyrA�1�E�f�7u季Q��i����!ZqcbV�I�F��Rj�����P
]�(�|�Ȃ�m(9@zh�C�� �c��Y�E��yjK�~p��;�Q����)��<���-����37���X��� G6�0��"�*\��0L���Äv��\��<w�*��^`�.�yˋl�J��Ϫ6�K:&�Q%Sc�K�/�g��GN\ t*U|�=�7���$)�[ �8�/ƑrZ�P&�6�F������Š�*����Ҝ��vA[�S������c�j�m�d&�@ (GN9�2�%��o�C�[�����Ha7H`b�t�����ψ��q�DO�r�����
��o[��=� s���?y�%?$���yF���d�.<T)=.N��p��v�6�Ecݶ6h��$��c9|��K5&Ɣ�k�Ds��W���e�,s&�ApA�Z��*b�G{(����΃�]U�{{Ws��An�����Vc�[���t%���V7W*XqJ�V�%-����[��=�3}���!'n���x*�Ã��-��AT�~�f�\K��f ~�Ų �p�3!.�n��d���~������B 'Q硛y�;�=�?.���EۘEi���gն.8�D0��z �p����A|�17�"~���H}��*;���Ѳ��j�����,�<tI��'�	&N�q�evóI����${q���\���7Q����r��y��Ra9@�`P:ǼO��2ĝ)���o���}�Y4���<�q��C����-�2[4����%�����6�K���$��Ɣ V;N	���AN���s c��Z� K�z�7x�}������<��O�Hx��}w������7͎+h�}��_�^��A_op��ǌ��'{��P:��6�r�n�@�`8��+��N˫���g����#SC��0;<̏R@
\ղ��Q8�Nu�cr\^#@u=���c
m)8�D`қ�����3(����������)v���5�z����TGN�����y�|[H��R �����_��U�P�-h�|�@7�r�b�憗~_�a�� �&3������MG�
8-0�c����"^L���_}Y�r�X	��#%b���_KԫR��]��矴X��9�ʭZYR-7;G�QJhp�#u�G��ԣ1���e3��`�
��z�2p�z�\t������� ��q�%��?"�7����Z�s)���u��N��n��z��dגU��\��v)����=�|��@�I��s�*�(�x�J������Ռ��ՖT`�7�!p1u�� ݜ9:� ގ ��xL��׽Wu�;u���X,���I��O��F0�	�/02�5ɫ�z'P?#��OC�/#?��Pל8Q$j����F:�����L��Bj�0����3/�Ltgg��>�1^��R�����,f�'�:ߴ/O-���x+��+�@*�ܮ�kO��`=�`��&T��k����2�Y���3�çˢ�O"鉍q2�n�SI��G�R��� �J�Y��tMF$�����dB,h��#�z��H�\C�L��Y?�T��6S��z�O<wI�aA��D������={>ڢ�Hx�# ��9�����#���8>�j1�3FI�5��!�N�<߰�g*��ka����Л����b���J�D��2M�~��s������~W��� ��AQE�a��b����Ǘh��.�U����&·��񛺑���i2�,���MЂ���!��j�w�-�J�q.�o}O�қ�n�|��,ܨn̷���L���/��� ��]h�<�a��@j��.&n�D���Hh:I޸�� ��m��Q��"8>*r�ħ ��Rޥ�rѿk����6=D�>�%�P5��p�em�|--����5��N E�r5���W���3S�^5�<����}� S���l��Z.|�s����4�ʥ	:�.�ݿE/z��D�w���P�n�^�Ȱ��
:xl�!D�59��n$��uA������V5��W�7��)�w�;.	��Ā���u�J����t~z�a�Q:1P/�aG��ت�7PI���sJ�zL��Цb|ʱ��l�*�$,>�p9zb@��rF�ӱё1,4�?'@)>����%P�Q��k�r+5���"t�t7�.K���Q����@'��*kJv^�u��jqTv����|MH����7����*o��&]�<>��<����*4ܭ݋<��
������t>��ԓ��I�5~�U8����z	Q\)�:Q��8ˑ?:�/
8��sU�*�z�����0�ߑ-�z�.��F��O�	j��s������6�{�+K	�_�´��;����˩��t�Na�{��LB\jb�H����9>��<-0�����_.o����"М��=V+�}���l</��Q�2N�|��o�,T?4!7%|I�%����l���وI�tJ�- �ɓx�		��䔌Y�CQ���ͅ�Gj%L�ۗX�gn�t�O�Rكm7X����\��k��qĞ�ۯ��C�6�A�!o	T$8u�N�3"G6�ϣ�,H>����<�e�C��{��i0<�,�Hw $���}/h��_�LVEЋ��T��T���K�i��i�͐>t���f�t�u�W:'Ϡ�9m�)>���Q�-x�*H��E�s�M>�j�����#x���.��5 ا��LZ^m��p*�Ff#�G�o�R�fl'�{ڐ
F��)#�f%⻾G��k&��&u�~Li��kX��q�;f��P+�B��,��#Zq�H��&Cc�8!��7T��9�U���ZCF��]}���ѩ���!5�mF����.CqV���{�j\ګ���ΰ�휞vIo�
	���7"󅢚v�����܈��?W��@�B��#H��q��D�C�_��, ��"��/�LoaY�UNjG��g�ʛ�U��ʊ��e�F,c]�C�6�k���� �K㤺�����2�p����)0o(�]�{��ݯ�jI��M��¦n���~�zAV�K�*��f!7����e�j�������Pϥ�-���=���[?%�tG��+��f֓f��ļ�"y3Λ��������x���'�x��+%�#��/!tq�?E}}l]� �Mz��,:��
K�S�bf������d�1��"!(��d�C$��<����'�k�!X�
�T�$�h��΁��(]vl1<�0����tO�<R,-|��U�^K�^��P`������`�(H����o	��E8z싪~6T�w�iJ��)FסK'�p���F���Q�Yr��}6�9I��<8t�9�ۜ<��ł4P�{��`��~zNr?-Ok���EH9�~ҩ��|��>��O�=���PD� GíN6pU��0�	���`��Ѹ.`6=����7�J�wz��̰�������{�$��� �;|��6�uN$��R�$JƢ����V�����[�W>ҕ4y�`��q̼�[�:�F�I]ԧW�����I	'��a9�5�$>����T�fl��P.Դ��k�ܪQ��z��ZbOQi4�#�c��|J| Kr>
VO��}�(��OɺN�`i����K�Ӽ՛�ɠ4r�����$x:c�nNi�;��E+�&�܃~�X��{@%�;��G��#�@���.����yR��V�Okiu�Q�L�
% l�א�*[+\W��ߊ7T�%%�j����H��&�o3y�G��� �OAq�j:��i�Q�u�%�����_C"W&�ZM&�Z���YA�������j3���f��c�'���=f_z��GX/��gm�{��FW��#����c	 ��ū�\CS���J�_�F��Д�~�x���Jp�5�-|˳n�.ȃ{�u�<(�2AW)]
��Q-h,'�q�_�4�Gα;�X�D:W��lD��D�E@���p_�ܺ.�9��	��c�v���!������PB
N�/��KI�����7-+6j8�E#�`�]Umkϊ���iL�nY��Ht��4��R�(f�`8{�eʣ*�wB���LH'��*�Ә25}�t#�J�����e{��^Br�Ž}	*�7"`�`cVk"��"`��6aɨ|��Bǌ\����+�+_�g���#@�SY1ţ��ݎ��fK*��n~��?C,�m7KW���>�^+�"nQ���v��4e�фD�*��5��1]� =�U� M渳�ޡ��K	�n=Y6����^YJD&
`�;��Q�sw(?sN4�0N1%\+�4oV��c���%��|y�΀��S 5��ޢ��)� ��?�5^3�Ƞ���g�|W�2��lZ��
�Z���1'hX��E�Ѵ��"U�����E,����rBq��0����֟������[!6`��R;��z��!�/�����*`^;��w'h��Ld"�A�R#!E�
܆��|�stQ��MoD�i�T^������k��'q#��+
M�&�Z/��tI:�3(�h>�d�O���\�4m�𲎚pl�4�>s ��0�;�l� V��7*RT�B��Y �d�2ގ3� WM����[jL�s�C�v윜�o	������U�(j��%d�N=/b�����:o�	��T�ʊȊ,Hg�aR	�Ǝ�J�B��Q?o>�>;��9�D�L݋F�K��E����<���>nQN��?R��^r��2�x��xL�+��-�#�ۻK6TrJж<ڌ:S�&�p�1<Ҁ����&p���T��Ybы)A܈L��co��BjO�xa)0M���=Jլ�~�5�N��L�NNn�fG�b��46�{ $ ��`9�I��'Pn��i�-�i~&�t���U9�!0���k;2�ߋt�Ak�.�	�,����� ���x�Z��4�}� �e2�-�'��0�lۘ˗�:�Qt"=���>�LSq9ښw�)�QsGPV��C6sb�����`��K��2���L2�j�/�W��3��xf���1[{O��d�X^��$��#V�8��h�����q!ܪx�֜�!��F���t(A�q+�{�X\G�y��Mjs��}��]�o����#��O���#<2Rb�ð/(�1r��7&	�O!��x����:�,��������k��tJ릙�(]pz|%ƚ�����'t��C����i%�O�鉶эhh�h��7�G��$�6�=�ⴲ�׶��R��%����=r0�
��300��i��$i�x�:p;�{���Ƙ���EG?vl�����WT�d!y��ɝ�1b:�4Y9�Ҥ����4�\q�L�4�� -�l	o���{��ώ�5r���=R��)�T8_��9L
+n&=b()5�LIR��J���1H����q����p2����J�

M�����G����ѩ��z��`�|߽q���`x:}�FJY_T>,SԜ E�|3�Bs?�s'ҡ\=���{�R+���G�@��Aȴ��L��W]�G��Tik8�]��o�G�u��LM#��W-��@�}���WT���j���і�l�"24�^�\�K*%��ŶʏK��8}�-���~hxQH�LY��<e�v�N S��4��� ��j۸�s��98�˝�E��LtiR���W�j2zh>��:�D��1��Lx}�lm +�i�DV�@�6����69=~��Hq�P��T���Pʘ*�>OU��]�:������28�FU�͜	�G��<nL�{�%W����&G�9��
�y�L3���>���7��aKI	���ɓm�Ucw�K˲z�j����@��!ꀉ���灡�7��`�UIz�<_�ޞ5��O�E�/~��>�n.�2�.�?���������q��*��a��ˁ�0CV�s�|k
.�
�ː`</V������[j��8���r��D�D��)_��]�e��d��r\Ư�"[��8�K���r�K�~�O��X��x�}�
�� #�)�m^}���f.��Z&�D�����"`����ˠ��n�d �W���7��M:*�.�9 �q��q�p�36-LܪBL#���j��(O�MV����~{����>�]}E q] �U�g�$椺$����y���=�=
5b�X�_amu��Em�ѹek�B�%g��W���g���ڡ2��札1ϡ��Τ�k9y�2�&M��%n��y���RPʣ�D��?9it]�H�N�sT�E�4��Ý�k��\/:?���v�')7;��\���xC�n�V��#���Ҙ����Mk11{�/��E�W�����v@=��+b����#SyH/�fy��C�=-
K�ك\R
	������lҭ���_ˋQ���S!3�X[P�j�9	��,��Oϻ�g8� $��� YPs"�]���P��Er�'�`��T�禶�$��a���R�Gn�Zڂo�>��%�s���h�g!��B4���}&��&;c�e{(����H�^_u񼁡��U����Ůȑ�=�t��� 2��������z�B{��7N������;���Y�$he�A��K'�t��`}G	#�����9�u/G��u+�J�]=��XU�G�Y6 ���!]{�q�o'._�@��ym��f�9	���y���7<���Ť��}t��l��x���zO{�o�K��l���1��2l�E/Y���ʲ��'SZ��+*ĂH��J\19�ڲ�A�?��� �,8nZ���{hq̕��(a�@�KS5��~�H�u�$i�H^L����8@A�}�����:aqJ�_ރE����������W�a�ܨe�C����<�U����\�Z��[M��#�`�F C�����I��Tg��������|ځ����	�i+�+ê�R�uLR�]�-t���,�����-�9��+1Z�<�N1�C�.�x�ۙ����|���!�y��/LP�"h:3�qqMU��-$e`̏gF�_''����4��M�l���X�)�f�غ��![1���l�]�1AGQ�ዔz�7��n�������s�z�C�L��b0��y �iK�$]�tE����w�k�u���K�m$s�晢o!���\̋hI�{6ף˷���G�F��ĳ���bl[`>q�����3��I���6WV*���+g��0K���9�D/��[ZQ�r'n�27��\%���3���Cۑg�nD����xB�B璱l�Z�B���-���阻���l<,cx��D_\R���]�n�W:��BD+�]������)U����^}�����-0E�ۙ{\�\������hT,��s3={�K�K3���<���MZA<�ȡ��@��"s��1�m�m�?��){}
�>���0Ӹ��n�y��O݂��#�����f'ĭ棆�pm3�:Q ���J�k����X�����Z̮�0e����v���<��}�^4J�V��<ג5_(�B�u� M�w���Gؑ�����h#���&��uq?�p�55Erl߁�sw�w1�{g�mȎ�f��c�0�b��k�C�Ͷ-4}�CI�������04�� ���N�~��it �K�2=8�+��N't�(�;�uP�ᬥ1h�Q���*4P�y��hGOs3�����D���
H`|W�[�v �tX��_;��Jma~�f�,�����{����g޿Uʥ�5(���@�b ��0�'���K�!/�@�IߊD�<@��|�.�&�cn@�ϝ�`u�����J{3yh�Q�4��)���������4q��]"`f8�b6�H��t�x�e��m��3�,�ctM\�x���b��j�*���F�Ӊ����ۉ��^�d��f`7&���=t��HPr��˝��E��76���!(7W���������*j�^�ek���MG�A���{>�YzR�̥�%�^��[&��Ǖ�h�M5�?�:s��m_�6��ԋ�P=�ox5���-�(��V��?_A���e��4�b������+C"B���������d�&�-��쳯(A�I�� ��$M`��X@�ïײnqs���bB���!�e+�d��K�,w"��B���e
oN��LX�~�qb�p��U>��j�/�x�� �)���ų�Y�s��.m�+W~�E��
f��7^�04���f�@������9?��Ͼy��{X=ed
ns�P�MN�R&*��wi�ON��9��o�8��.����W�W�"�"��B��.
���E����s�L�$h+���2�� C�C�q�05������L �k���ˆ 8��������
���ij|�}�?���y�s��IK�%CC�������ᅄڗ�����/Ҡ�XM��  V�y�,h&�)���	u�93��<�iF�	�;[�Z!�,rmw�	�Ŕ��Da��n-�\����[�����,�b���ԭ�cd9"�j��,�׈Ǡr��a�c^���Y�=h���Ej���4-�/��ӑt�؏Y�ً�຅�E�U<z&����U��uۯ�=�f�,�p#`�/����z���|xr��8��Ҽ�����
,UM_�ǭ������렼4��Kn�8����G��w�n��8C$�cTK$1�n�X��z���a��]��#)���(W	,)�=UG4e��s̍"�s����Uҳ'�S�_Ɲ�C.���J"3��s\���\u=W�u��	p��b��R*�1�n�u�Qu��`2��]�"�ߴyByafӲ����V�>ꓛ��o�,�A��2;�?1��Y�2��̓Cx������|Y@oe���Rh�~-�LNp�J���V�!��eAOu���_�V޾(��W@�*8*3N�� L>%Z�CU%|�wO
�� �݁��{��@��ANN���b~Y�]��A�cp}��XD�!��y\c���>��yKx�����0�H6��wj��S~xtK��Џ��xP+Ğ��;'�p/���+�o�4w�L�'��6o �P�ٌ��Ol��춍�@͋�O[�i#\��ٔL�&6
���>��t�eＧH=.OJ���RF�C�V9x�b�z�D����z�p!gn�(�#+��d�RS��Zp�g7��
�2�K��Y���]�����y�[٤��~d���P�nEcγ����d��Wdd��~د�*$��]m�x�Z����]+�z�r��6 .9��'Q(�+���N�M��<I�p�Tr����b�u�%�j�=�{��u���� t'|��B��ɲ�W�B��>�Mu����%�JZA���*�dI�?ϊ��|�A��� �~�;u�wS��6lK��"�2w!���0w!�sm��1�j"_����а���}�uH�گ�a�͔�'�^�58-X�L�b��~����gб7��wW9��K��A8�$��ɾy6�Du#px�ք:�T�b]n����oVnS�x��Z�Z�������}��]#�Ȣ�����o��T
��e�GS C�1�(e;5�Z#��.	�.nSWqn�$�=��y
�9����J��Q'hӶ��4�,۹D��L�&���.��zӒ������B���PU��G���j%����D��n��/:jÔ������ݮ����[K]�L<`+�;C��3>lݶ�'f��ȕv,���"}믚�YC�j���cC>03'����p:o�IJ�<{]x_W5Z�0'P"�;.dezEx���H��ON�u���j�i0ݛ�B��L����lt�ER�[L���52�j8�25���..�h!�`7*$�0�����}ݔޅ|t<��ѤDbuX��K�G��h���{%�@�f��ij7����:8;D���m������5�\�j��/�����^�����g_�c���QJ�	�X�&�I�Al*v}%��r9���g���\ �	��x�)�!O�R���U�-�|j�n��&��\³��H?�H!J�!�E���V
�7�N#����DDq�_�_�U6�>��и��Hd��l��~�a��`W,(>�Y\"�z��Z~�����_$��M��^9]:�F��*zg�1��ԑ^��HU� }_���F����a[��#�%�o��F�NA��CB�2*�"��*y�	�\��d4M�G\��B�2:��lδ^iaڿ���;��p���됣CK�q�Ԓ�_����Sag����*+�X��3o�1�t��GPʐȦb�7rp�M�  =e\ Q���Mbt�B(�T]�m�	\@,���SJ������$pJ���'� ԧO��)r�1�~Q4�(M����<F���Y7�w��&:���e��I�׽�H�w�w�j�� �8��1Ќ��.>![���Mܢ~e1^M�=1x&�s�MG�+�ͨ�..9HY�r{,޶`(3i]�C_y�j��A�`4`�%�`������*c��kͲ�uT�������7^�:M�7k������ƕ��\�J� yx�U]}��˱h�R�T�}9�.��L���]aS����J�k �3Z4b¤����_A#-��ݮ�+�c :�&q�O��'ˉ��^��]p�N{@	�Dp>� ���I�烵DY�� �;7�,�.5�5Q��U�~?�z�/��r����^�ԍ���"N=�|M�uuE$��5�rySh�'�_d�zGF(e{Zz9�/`���$o2×X^��%�� P{��  ������-�	YIl���	�Q'��9f�����D�%8?G�u����&@!-ʈ��N�XB�j9=	���gM/"�:�g�!�'N��(ۍ����0F�}�m���V�Aݒ5E ȷ���\�:@~������e���I�۸T�n�hX�E>ӠA���?�Z\A�?�!�m�J#�`{O4u����S�v�_?����?/3!�fdg�j���a��r���ԥs��}f��+�0�[Q�5*�FY�$�#au*��r��)��������Q���2���[= ��dlv# �sG!��ʥ,}�:��9�p���	�+R���@�J��W_._XFB��ӛ�ڎ-�nԫ��s�!�[-��&�Ƃ���ݳ�C�ç��Zd�r��Y�&�9UcT��Md	j�A�	:q���2�̫?��T%�Dd�܈�ׇ5l���آ$�Y<e���I��
�w(�����.�'�m��¨�<�����a9(ځ姎��lt�ŚA}=ʹ`AX�L�z�X)�/_0->��QĖ������"���	s2lzl$[rN-ɿ}�ל-P]+�x��Og��1
bV��� ��N��oZ�w�uY������7���|���Xj��#̨���7uz�*x!?D|�d�ji�Q��P�&۔ ��h�rV��;���e�U�z�n�Ӓ׉��a �gt$� I�0����c�!��� He���>l����Ұ=��T��?���>����[�͠Y�n�x^8��pP4��� C��f�!����6�D��(�m)	���r}��)��)��~_���`��6���V�n�?o3Qy>ef�� ���­GH��,���I5ZC�U$LG��Ǵ��/P�G%��)Ơ�D2��RS���.8U3�ޒp��eyH5a��N'����������l!��Z�B$�.�x�7�`�p��&�y�+j�,%D��C8~��$ce�фϼ/k.շ9E��C���PpU/��e�:�oTN�!F���f�&��bc�A��3$���a��H��	b���䩷�-�&�bh����0i���#��� ��g�#>�]��yK����Ȭ��N��2f�,��|�2�_LZ3װ�*���b���eR���=��'�7�z��9s��y��g�>�~d��z������c@�Xd0�����E��}ͺEnd��I5��.�B��x�(��nyW�̝�q��V�ܔ&o׿і!m_%�,����68��)X��u�@�����/YNmv���(K�0)�.t�/.���
񳢗C��WP�J��rv�Z�N�ڬӛ��+q�K�0��+�`���D
i�h��ѵ9��v�+�^���g������d8`�q@
v�~=�y��o�<L!b��{GŠ�挑�V��h��q ���O���מ��S���Y�����5~�O�U��^-A�Uq��oA[1p8�*��?��	��@pi�־IC������h���$�����׻��tR���DK F�h����4�c����_Ej�c�u�E�h#���t�g����D.Km=��[+
b5w�����U��8G�D����3�>)���k>���0D�i~��L�qT���8Z*n{�	�� +�C���y9��@s�i�L4x&}0�x�o9�1��1��2VM�!��\�f)t�A"�y2b�*cK�hc8E}�±%�`���O�'����qǀq	�"4�X��M�����l>���C�J�#������;OS���P�>��4{2�
���-�y���\����}� ^-����#�a�Ŋv%ѳ�s��}-�!˸g��d�8H�ı��T��ࡥ���)����xC,�WV�Pq��|ҟ��92��
 N��(�0J����˞����x��إ	Rך�dC��y�%B΄US���+5u�{��ՌkBP*A�� �Bw�����]�=o�M"�;Ff�&F����w۵��Qh���6:&�ƮKc����ݗ�uP�+9���-!��/H�EK��?��#�����)I9���&l;�E��Y��������n��?�ף��s#���`k	d�'�f��Ɲ��]׫&Ov�Yڲ�n�m�e!|�E������ V�kI�����:mXz�q<2㽓��`4e�^�O�������Ku�na�4�>�菰V������Ƈ=�E�����t�i�� 4z��&����j�1���`]�g
*�w�bGJ���iM m��Sz��΍ۛ���2!����:21�u� ����g c��I3�Z��0�����r�j�|�L��p6�{� �(u��#<���Od�s���U�Y���݋ܡG�x���X�����A��j��I�J���X֛��1�t��nf6���ސ�o�~��2с<`��P��w���\�з�﹄�]� ]��E���:[l�!�Q���$�]����}�����(�-�~�L�g?O�tb��C��d��������!E���A���o��5���St�9���8�Mc�.aތ:8rxij!����I����{�	̇�\q���W��Ƀx�!�Ȓ���)��!<è$T��b۱�eô���t�o�\���Ї� gM�tO�o��f��Gٳ9��OT����CP6�Z@����Va}H��t)����SFQ%��� z�ӆK	��S�����&�Y�oV��6���OOaܞ$[~��Y��(0�O�����O��o�=2}�f-��RHp��I�tn-���x�"�ÈͦkyC��a]�x�+"�H�y�s,!0�ٞ��p���л�=����R~b�� ��?�$��b��EǸ5���+L�U���F�&~��I� #�@3h�9��m7,�4o��1z��&9)J��ү�:͇�ۊ�o:�}�$Y�2���;�3�7��&��S�J��E@�Zlh-�]�Aw�2:4u�3�K�3l�Y#m�	�xP u�$���V�g��}�.c�z�1�0����J#�A��=�b�ADz@'t|�]�6׃�[/�����}�`��r*�a�H6}Hii
k�(Mzm=��c�R�b�;�(_O�Hcc�%E���0��<t�]v� !%�Y��S-/<,��GL�SH$ԑ(��P���c��w���j���4�ef��Bv؉���lX����摲+�������	�Ρ]b�s��?�dB�v��Y�;�M2�-I�G޶���_7'������������V��r�ʷ�[9�I�ҳ�9i��Y='f�P3�U:�� ��mQC)�r�V	G��;'=��H���+6bI�2u�r�u��-?���M?��I}<����s���߫��uLfý=fF��fD�~����0[A�I.<~(��d�8�="��j��T�+��Y�X���^�?0��(S�X;`�XP�ӈ2��̯5bj���C�q�;�0(�o'�3�B��]�[S�^j�B�k� *J`Q�tъ�X8i��c�.O�7����_l1T4L�K��ᅣ�a����>�SuAl����O(�S��Z�t�'5���.��߿�_g)�d�驊+��p��(�A�P�������!+lk��=q���p�֖�`�`�m��e�h+�^�l��j��l�0�y+��\pS b������Χ|�BXؒ��y���O�4�HP�2UX����~�Cr����&u��Fޚ��{<A�&�|*i������d�Z)�N4ꄲZ��r���3L�T��wZW� W�����"g�}Cd~���MeP)u�n�d�UM�� ,�K'�B2,� ���2P@uR>\򃌚���������g��������]�~��E�=æ�7^%K�pC�|�7Y]�t��&y�s./t�"��x���Ȱ�<���!to��yQx��G�vN�]��LEY���oT氄D�j���m�4 ��zW�Vޙ.m��O_��O"΢������?��[@�����#��8w{7�<]�P�L5�%������n?��8�5apT��4w�k3z�䒷Т�[��4�krK��w:b��i��P��rcڍ"?�ac�%�Oհ��y�jE+�xY=Z^D����`�����qFC_�0��h����c*���{3b�;"rާu�"ֱ��׺��ό¤6~�E���΂�E�(���1B&�Z.Z`c�+��w�ѫ�����/A��W�DL�p� ��߀��P5�q8������צû����`u�~S\"7�O��q��g$N��aLF�����.��r�Z��Y%T��3�� N�L�y7C�R���g���+f��A�Y�?�i�񎁚���O���ߊ0~���<P2�X0_�X�����f���du�tz�?1���#�<��ن�پ_Xn�*�]>���㉔#��Z�ԯ�;N"	\(Lf^ 5����u�� ���5��y��|Sj���摩���A�z%YK=	��½�Ii��+�ZLە�咳D'���b��=x�b��D�v�M˖@M<}� {:v�9D}U�%����'gg����ǜ70�w��s�S�~��k��׮j��%��M|C<�OF�o�6^'�C���>$p�H�{*_Q+�x#��C�j46�p���*�K}�R;ՈoK^���	{��bSIu��6�UK���<8��;?�`���A�I#��S�Ծ���AR&PJ�U������ٷ��7�é�F���W��5�2\9vОR�o�:JKȂ��1�j����:��Q� G��
G���lS
�c��i9��M:B$��S
���R�jF���k������Ҍ�i<�'�k�o@��z��y��K�.z���C,�C���e�\�?�`�z�[G��o�W�n�r���@���|�I�HY�)	��p�j`Wl`�<�d�fz��{qI��F��T��2f�f�+�&9��KO$����z���x�l�>#�Z�/G�\�X�����rD��.W�+b�1{{
%g����,�I`���X�
 ����%�����ߚV������3P�u��6A�^}P!K�̚WY�m��&�K�A;C��g�%���e�w�[�s9�x���盩�J.����)n��Z��`9
Aؚ���ٻ��IڑZZo"i�t��W�6�`E�$��Ȅ������t�ɩ�C�Ga�1���QG�N�:/7sN0�G|�A�"G<|g;kMa��_V�h�ܢ�??F|�eC�L�'8�&n�)�Ҕ�[4f������k"�P�,��]��ޙ��Fc�6e����Mw��vxܢ���N�MIΥ�7J�YH��iH�8��x��� ���� ��?ry8M&O�7\�~��}3��-n�F����Y����8�"�h�.����EO�a�Z��(���7e���K/%�GDʖS���h��-S>��c��S�(
��?r�3��X�JK����f�����'��.�EQ!*�C���s���f�`(���Ѫd�:�e/�(��@�g��<�ڪF�A���]�������OGcW����3�߭��Β�輙BH-��羷�
_Gԛ~�[�f6�1Y��c��;�}�l>j�Ӌ;�5j���8\$�F��k�6[$V����J}�� eF�����8�,���pņ����x,+����P�����<[�$ ��զ��$���ȿ�ߋ��R%��_�a����!�Z!ƪX��t�/�S]����m��w՛��N�2��h��OI��sB?V��v����]J:4Y��"']��}̣oI�|�M�:�e�x��Gc�J�S��$��)s�I��XZl�.�&mW.��4�C�Ѝ�Y���$G�p��޻(�z��'_j���QV�V��'�����֔R�%Q��5)]4i�ze����:�2��S�b	�S"�6�n��m2��~��"{��b�E����
��m���iZm/��J�;o���$F���7H��ȓ�7�BE�墨Rt�IDC֏iȃU��w u��j�����?b�\`�I�ȋ��c)��]�$~��2��m���1����O4��Z��e�~�M*v�y<*�H$����dC�S���%k\,"��S!m�ݎ�S>kq=Ca{����)��7n��>�۾�`�a�6�dz[�r>&5�U�y�%sq��
��Ģ�:�1�R�^���G9�ߌY4ֹ��5[Z�<��g+9/���������m�+ɾP��7K��vc�z�WO��m'�J�/�l��;��5W&m>?��_.�l4��$�N���=X�v�u��؁���q.f�Z0U�m��VB�w~l��(+�YOh W��3p�����+]r��k_i�M�[if�Ɂ�V�,�����o_a���lnLF��DԊx�TW+�⋹c �����/�e��`<7v^7X/�d�6��f�[�kn�#k�H֦�Ԝ��kI/sdW��0��5��4vp�t����+���qRy��@���KB�
3K�럋u]��`!:��'�UY#��dY�-��K�'gd-*��ݹ#����Y��/� ��TWD�\f�������B�<�� �zV��êh�4; �&���{63ɥ葞�k������,��̘�h��^C�aO��f	��q�0��~�S�pj/P�
��ʿ�V�m�Z
�3�T��uǑ��o�(�&=�"�"<�9�⼂�z�dڿ���x�x����0��<����(*)~<-F������ox[ǋ�FiNf!ᒼ+�k�����h��A�ynl?��\]���3��>˧O�h����2�UU�5j1������U��N���j�����ȡůk����E�+]}�)x:dp�8��ϥ0�`��Q���aM��G��'Q|llU�ź�=2�!Ԥ�/��u� �bc�*�8�$@ ᛛv�w��X�3~�;��)��@�yIٓ�R� �7��3�R;���fַ����*=��>?�����j�#E�P.�շW�t��S<散c�=�~w,��P�A䜥��Ow�f�_`��4���=�߹�+�9�;-����ᶑ�k�ޭ]S�yGY��W�r�����p����]	6���V嚊H�|1��y�h�(�`�&ASgy:ɇp�Dy�c����3m�%��0����6���1�X(���-��R��������z�N�iac��E%�YE�[�R}�|y��^.���ZS�}!s��6��)M�ڨx���g�'��J��C�l�!r�/P}�ۃn�x�~貅��?��8����W:��P8#P x���Z�����'@Y&�� K���\S���kӝn��+<F�F�=s�Z��ұ�\Cv�f�^���@��
��R��>�F=4��UV;+���
 U:��|��UJ�/q���g��d�.�P�I�����7�$>��]�~���%�ut\���HT�Y7�Z0�$?e[�ԫ��Ϛ7:���,�F��#G7��lv#n'�=��该��%a#�j-*�|+���s\��Лd��!��=t/c}�NE��\��j��d49�V�;3�/�0�V+��;������/��Ε����*�}��$Q�e��F�C(��켡=_���H��h$�6Sr@���{s��3�D��D��;�9j�'���ū������~w	���F��ډ�r&}jA=�'
N8��R@��~|��ڽ�ӆ�eJ���A7� ���h�K@���"���=%���~տ�JZ~��zDM��\���UD֔Qe�\�/}�uuâ]7�����wA򊓹=�|���[�e���J$����;_�ף>�w:��M�������n��t.%{��M#�h�\\9�z����LA���A>�=� �2Ǵ�n6R�8}dTl��+�7&�=0��MB�Cu��fR0B[GLDǔ����lP�a9F ���{6�9υ�K%����C���,9�c�\v���z~������iu�#F;�hq�x�GԶt�R4�2��5� 
���Z��i�����	M��D��v�� p��}6��x5O�2�� 71���3�;*�X�X��>�:e��-m�§��_k�з���$?�^��#o���}n��w���84�N���e��e�򁎑�!��	
9r������
�5#��xx+C|��-�k���,��9`s�	x�ހ��w��G<��7o�U-`�\ݱ���v0��p�)�a/O�t^��+U��=14�����k6����qb,zDsv���!�l4t���p$F2�F��Ax!��8G��(p�=i��i��Q�W�3���Jۺ�Q�L-���+���K��w�����gA(�V�EN��
#����=���m��5�5W$3;�]\[���;5|O���v=�d�Mץ%d<P#�Ka.��L�X<oX���2��2�Wh��y$�ƈ�5�l[�k;e��yV������x�#��"�������@oV��nn���CuլZʥ�]�k���'�.��� l�λ|���^S�(ʩ���D���c�_�
�ˣ���)��Ϳ��q(�Q����e;:Nx lg��UY癃_iyb����Nb�u1�j�^��~(�%��q���x^Bs�e�%��UR=\�_~8)d�a5B���
�ge�mj��by��XAq��&��w�e�����Q궢ה>o�cok�>$p+�x��ҙ���؛�Yj6����z]�4\�LB��T2�F)u���2�@�@:��b��9aUٿWw�����w6L���ڣ2cX����+�p�B�UO���j.��6^[�gC����n��Y·�G�sHA�,(�p]�����|��`�)DK�a���C�p@]T����׾n_my'J+U;}�qc�w2�4t�o�	��Io��H�Z���X�= ��=� ��w�#j?3�%F����K��^��"��=YR
nn�d�� u|�y$�/�Z�MM�+��z"E>x���o���Df0њ=��4O�m����4f���i�~>�9�n�uv��CY��T��H��Ow�;f��a>��TB��pD��"|m�6���B�
b7��=U�_���9�ہB��E�W\p�����GJ��3,+E}c-�͗�n,�<�~���v��6�fO��0�<cs��D�2uh��H$/-�����|�a)�ߢ��� ��I�n)�Q7�c;�Ue�za�آ֯���w��u��b-�G���B�O�4�{(�^08�6k۹�X������MN+��"�*J�t������3��˹��A�HvTɯ���p.(���^�0��U3��c�c���\�5��r&�-�>��������m�f3�s���WH5�c���j���Т�q�����<{�w@CM�B;������.�U�RckM�ٱ<�?��(�����J��T�C��]A�%�.E�D,C3���_B/-f��7y���o7iz��mraEe1��^�^Ǥ���%��|���)�ְ;�X0~/z*��d��ll;���5��3�{6�Ò�0��d��7�,LKO�E=����'��M�)6y�3$�\zb�{G���KvΩ�loذ෤��^�N��񩳮���I�Oќo�U}�%��dHt̷t4L��?��$|�iL�W�!N����n,%���ߒ�f�&��Cď$磑>��9e�v��p0j��n������T�؏5�7B}c$�F%v�ǒa�s0�D�����-cUT�M��%xd.zZ9�`��c5̏�꺍���kh��O���4��o�I=�)�V�Va�T�N1�@2�u)O��ڒ'�V/-�@��n���o�kI�Ϯ��'�$9��G�j�I��x{��lrwg�<� ���0�i^�G=�򢰓Z��$w�GU��塼S§�JpWv%nP�Agt����Bs� d��nko��u-�Y�r��w%��0��)fN��i�d��^YY�~6*�BK��S�>�,Sk��h�DRI�bv���������ߎg�۬S�=��T�Uv����\���jK{��j��N<i�tR�G4Ak����2����48�R�a�E��E���H"g�1��[V%S�ʚ��m�~����=�eO�&�t���W�p6��}3�G�Wnf��L�/L�Q Ϳ�|'ΡI
���~(j�8�1��zA[1��Ņ�<��%�؎��O_�z����b������,�lw�H7b�c]l0?x�)�[���o�i�ʻ��_r�P�3��3�"|��+��Z\U4��!M,S��D�FR-�&ӂOf4���j��A����w�7\��;&3�ܧ��	_����͡6���rlE����L���U�b<{����
�;w�,O��Q�����3iTUL����(����^:�^��?���Y���Ts�׼TF)��]���8p��BѤ�pa+4Y���+zL��0���u��l\�[q�ڹ��H�oa#��k@�ݮJ�P�OuIҐ�P�9����)A'p$�DP�{Ԝ0l�:�?�����]��J�Ŧ�^ �I�S�O�Hw�i�s�n�)��_���kV�*%,(�����@�����C8�ܟ�Q�/��r�1�<�fEV�q�9=q����݁8ǔ�ʈ-�w�6*D L��p�P؄�E,��4����j3"�D⌑��HKpK�6����*�����t?�W剈�̛�V��M~uTԱ�\}�M!>U�]���xU���\�P�w�r�ɍ���EqZ�����V�Lb�;*˩��y���;@�d��[yVHF\�1��Ly�:T��������ᰱM-���d�w�,J�U����p�q����>�TBfG���Ί�Ƕ��g�#m..�EN@���ӻr{��]TwS�\�����a�$c�lb��Г�_p?�_����!_�±�L�5V��f���%�7��J���`E���`�?�c
6���-�}�x����1⾘!��!7��j����� AP����/>B}`*�B*�'ԒX���c�?j�'����l�'HK�B����je��|�}�$+�q�L���o ԯJD#��C�T�1=����rcM^��1�I�uq�e, ۺ�\(kAj4��gyV�P��x��I�e����1�:+�,&�N�r�V�{^�V`#�G���TΟ��\�?;�4�E��:�O��hH��%E�f��+�B0���Oߺ,���f0�˂s��=s���gճ�5�
����R���U[f��,�~�E ���q�"�3`��8�f��s"��p� 0V	"�� j�����3��Y�X4O.�BǮ��\���j�K��E���rX0�
�T��#B3E�h��x�"�
��]i�(�X��U>�m�	�v�s��YA��Qv�)k �.h�#=�0)o�i+�[m��{�gn�z<Ut8�Q`�*��
5�m�R�N��4�'��4�FK�)�A	3z~�D�/w �+��1�'�i}_��s �-D��A�tQ��7�|%H������y���%�բkn��)	�<�U�<Ú�r�(U���^�k��ń"j|r��\�����3���{+�_!֓���|�%���p�c��ד&�i�K��d)2������`���O��,�1<�ü�YO<��d3U��Mq�����]�E?��X<�Zf��ɫa�t��q���W��UФមu08��9�)��c���.hgZ���[��Ҩa@I6�뷖*�F]	�uȬ}�,�>��֎�ac��w�!1#.����5�X&�� _��y2���F����c�Q�n�M�U�ϔB���;r� ��Y�m�ab���Y��<	Ok뎈��-	��a5P��T@�[��Y�F�)vr�`c��C��6��,��!��<���*�S��L3'�q:�^8��E�b�цCuc@�DSu8U�������/�w�!���skMJ����Gx�&������\�9=������zӘ�z$���c��v>���G��&�!{�>�>���R��� ۶T��P�<$@m�V�\���ۆ̴ ��+}��Q��H��Ia�jT��g��\�2��r������k<�|��E���w[{��ykq��>x��t�m4��Zo7W����>j�/��CR�D�e�����z[�����!,�0���M[a�+�p��G*Zx[۶�?`fDB�\��NU����{��������hX�GM~��D��<�:H[F��-��O?��"�n'A���iL�����c	ޔ����/�^����v��.�Z{y7˘:�$]: �o���n_����"��i�7�p퀫���L��*�R�GO��t.a��&��
%(z��g��fn�����\�\	�yI[,��4�?{@��qf8�~��{Sك^h�7�
�e?~֬O��v^�o撋O�iI��;� ���?������W������kMY�Z�������YR8't���]����e�#�h��n0�s�ITR�s��s�3���˞�$�@7kzc�'�[ӡ�
\w���z�nFRsK[��g�Djh���a5"���gW�84����}��,� ��	��X�+����e9�(�_���%}$�U� W�v-�7�)�@�;G�2u�;3�O.�-�<���I����O���7�3=	���*�K R�q���.����a�a �WY�ᾴw�=2���	\�?Y��͇��/�l��^���<��
<�/���	��z)��O��p�p�zՖ�&$l�6��dP�i!Y=��@l�����J��=\F�%�pI.���q�q[�j$-DC���'�M�y�s]����ʨ�����и��z�u�ч��9�vM����5�����;���S��|E<���v2z�shCc֤MV*_�u���:�J����x��� �����G���^��H���n�3.M:�k_�e�)]R��LB?��;ԏ@C�����Y3��S��{F?���s#=3��ݧ>	�
�I�����s�mk-F�$�v��w\��j+Dv�{��[Nѵ�1�ǁ�#�X�*(p�������i51JwI^�|Ȫ^�5�&=����V^HJ�w.VU��{|�.f$T�2F�VQ�o�!n����z�8����^��v����0$�l��ӿ]�v �� `rxuG��ǪL�b�vd��ț��F@(V����4��W��� �'�i�n7`�B%�ح(6��F����o�*\�VIh����U]����Q�wM[����;��Z� �ɜZ[������JLA&�����B�v|��G�Á#�<\�K�Y)6�t���?Tʼ���JLRS4�x�	)��H~*UE�%��cޞa�B���T�[��+R�u_́M�U���m�j�Ʀ���Xd�������g�H���tr�7�e}���@�|���s��-��L��G3�vh��3t,M���HY�G��$�HS�E������d�>	��
���e�yVQ��<U�i%�ZX��{Ru���:�E\�����S*=W��]�V���%����Ae���B&�SSr@����6�u���X]�e�oΒ�ּ�
2/c��[詺�h�^I������q��A�eii���t��oM!�K��%��3�j.�I�A�[y�^�^d�S2��n'�>�jb�G�Gk}+�F�lm\�?n&��mט��N��6
���r�Oԟ@V�����s�`���ï��Շ���������j�s�"�Bi���c�;��v�JҐ?N��Q�<��DO�j��2�8tQ��SQ�ѺE��9{U2�]�9����]��m5���=5/]��8=ґ���<�o�ѯO��J���V�PD'�ώS�:�H�i4���d��N���BϫiN�8Cꊷy�Y-=o�ucxd���h?���A��$X5̤X�:b�d��
��ܤr���/U��w\�qd�Y�f��iRL��~a�L��}v��/��g���(�m�-��%v��qgC�VAJ&0����l�2<�|l L�?yM����1�����ƭ���j}�6�����RYT~l��a��Xd0aZs������$*ƒx�q���3�^q��L,Z�(�*�I �50f�/%j��jY]�	�G^q[����4���:؏�)j5pߵ���G��o���w�a��_H�ND&5�[�s��Q�D�D��l��0�8y���"g]�.�� f�8{�6�'�=�A�9����˨���������u����6����{���@��GJeMi�Y�����&,��Z�����n�2�
Q�H@�)CUA��������L����{eҿ�����M��f��ܽ�/$1Q�ND�w��S9Wr�4�@���4	a��ǢI�:9�4{՘}�.�4�&G%�Y	ȈV���+�.�U�u2_>o�>$ِ	�R���������Y�.��%��.{_�DCt5<��J	�pl���m��qg�*<�Q�rE(��xR�����kS�}t|eXgft�]� ������"�"~��5W�U �1�5����Iz�:mj�K*�^8��ś�=b2n�lG�k���z�0�wi��*��ҳD;s讽E�ԃR�ĭ�*���%�(���]�:�E\�F}�6>m1]�X���&�?bG�9j�S\�����6Gz�ό��p�Ӣ����]c"\������1|��}�<�����B�Ub�����|*S>j�ws���s�秈Ɓ���42�A����������?�=�t�㕙���%�~a�%n][aZ=p��[�r O�h%p�u���M������s���O��ʐK���<m�S^�%$Z��� ��6���z5��Kʅ�M�^CxF���C�D�:M�[O;�M�!��a'e�T�p��Lˍz�
�K�O�i�A�!��Rh!I�x6��U	cnȈ|����M��1����k��6�v�s��f�j)������~��	B8rhV���ཉ;���h*�u����1��6�9��G�5�Һ���C�p��D�w��-1�t>�Ҕ�D�~q��|>֋g���n���f��'��&m<�2|�L�����8�8�R����ZTusQ���!g�!i�0&C����<�Y���'>�>{F�[�e��wjr�G���z�z]�KjLOο!b�L��/6�
���:�A����U�|��Sd���=?h2\aY���/�����4f������~�-����5X4�r%W0h�F�q3!�4�>��K�0˷M��lf�(2��B)8��eѬp��Z-#vFr����("���x�*�<�x� ��?����ajtҬ�t_?֒�.MJ��� ��jluv����Ɇ�㖎�F�*��p]�e�~w�-$��1�l�![S��Z��@$�"U��ձ�)fZ�D�=弁-��=5OqTň�u0b<������4ˬz;��A�y�����kř�.��%�Ԏ]L�μ Y�p����oԏ>$֔������|��!Ct��� UzԪR��z�`�2����Olgf�
,�ˇ��������@n�i�س�=pOAў��ޜ��;&N��<�l%D�N&5W����`yEMBȂ����˰��|sQl܃�8�0J�n34&iVկL�T���sd���,�7�8��c���k}����J����.�o��q�Q��0r�K𒑳��kNn��		�ӊ�L!M�t�c� 9���s��U�4�Ш�',�}gԜWx�����P	�B�QݓCc.�ӵ��5AK����Ox�7�Ҁ9�!sͶS5m
%3�nl�#ET���C�q>��/MYKh�������ң�⃀DV����WM�H~���׉��@���=���`h~u|s�)8��圇6G84%�֨�]�`>o�, ��������0.�>�a���;Q�q�7�bV:/E�( Z&�ELՅ��"&Q6i��l�En��|tR}H����ɐ��u�X�ҟ߬͹�'���?I��Lt)1��oB5���;N�xx&%xT2}��q9�Q��W�9չ_[cw0OBaf�"V[�٥��D3�N�f�&�f�k~*���|��U��PbZ[������m<��c3�����k����a��)��9�jr�:yN�S\���k��������V����\Y4T���czئ�ӧ3�e^]l��9��꫱mZ�A��n�������[����yn�/`)D(��j�5X>��2@�����N�� Ö�;���9�<���P��=�����|��l77��=$a,(�O��L��MN�MR�x�_�5.�:@�i,�nD<&`�+����O1n�����θ�iPn����Zc���8ra�e
���Ɵ�+���HD���f4��ͩ:Mf�scQ�(���K��Š�欠��ՃC%���^�*�6X���C�Z�d���������V�k@��I�9n��0�t�xԀ2>W��	����Hr�[����Ǭţu�[���l�3���rk`
Bk�T45��5h��������r:�xb�l�=|��bx��Fr01����/<�~5��F<��ˑ��wJ���ΉC��t�Te�=��V�Ex)�f@�\��O��yx0��dN���9��F(�z� �f��0J�3�/M閍��Y�5�
��ဍY���碦>�8x�v�/��v2WK�ן8�S�y���x�f,1`��8{������۠�`�Ǡ�)�{pʂ0H��r��}3C�����tE�AiR
�d��j�h6��ֲX|�cG���o'���&(g�ŻEl'�͗�Q�H�(��^T�����Q���U8:m_n�G���W� ��Uy���Y���o+Lu*ɐu���ޥ��3�e�d�/iU�2��n^FL?$҅��_��O�������A��̲E�GW��I���jBf����U��2A}�q�I��� ԁ*�ɕj��g��3/�#\?h��D���>�[Š�Z	�9��T�����;B�؃T��)��P�߻�;v�l�e�K +lĆ�|�Q���Mş�;��д��&t'g�Kd�q�*�����d��).,���&m(���Z0K��'�)M3�[�4��s���؏�sƶK�T�e��4���p[�6�>h��}�A�"���:Ɔ�������mJ�\�� ����!���b|v�;S���N<���?S_�0@�&�a�db(~93�{S<�;S���ǍKe�^R����o倄f��#�!����C��+����0$���i�{�V�C�u��ﭏDQ�����KY�JFFʫ0�c���e&�z��q/��w%4�}_�8Xy9����,�*eȇ�!�u�>Z(�)����	��@��ȇ�)M��޾����NxI�o�!ks<bv@��s�fb�t���,8�0`����c��V�]�����pu���3CA�}6h\ﶚ7�e�<��9f��.Q����c͈�f�����9/yh��<��=2�'t�D�L�,;�u!	Ny*�k:>T�@[5_�4S�N��e�Q�<�	�y�h�v���ǵ�wG˔��B�M@^dc�ԡ7����~<mVEB#��t���� Y��7&x��b75Lb��g�Mdp��R�9,��G��{�������e����l��9�Nd���o�˘M��c�H��Q*���N�u�4�g�:�.�{?70��@�vm#,��C7ڮ�5��	���X�ȫјҹK{[��ĭ�L��6����̊�=3RU�RZˏ15���<�=�w��r`|������L�k�J��LZh�<uJ��ydx�2����[����0LT�u��ɂ[K=~q ��Q4�O?���0Y_#E?�LK���rD$���}��}ٱ�6��X��8�_<ֽQ��`
���<��5o3��~����O����n�4_�j�Q9ѡ���B㳧��) _?�\�'eIy9�f�GdG�[b���-��h�t9�C�� �X��l�����m+�򃕰�dY���3�GG%��=���,�Rl'�h4��j�AB1�DW�΅B�\K��V�4;�~uT{P
$YGi_j\(��WÆ@{F/��M]���w�g��� ڰ�iXi�c��P��2�T�(I4��n7cޑg�:���K�ع�?��<r:�-�I�0J��"�R����`�O?� }�g�%z�&�]����-�&ጄ�Ur
���$��jRdoP��)06LD�$1� ��4��x�K�͏��%�BK��b���+���
C�A\3���
��*R�nP��}�b�l����`�s(��S����z/Uʮ[�ҡYyJ�HK�Q���S��~'�/g�g�28Ж�"`(�;�p���:�r��
Ҫ��J� �u��zS�#ҘS���ǣ���K8��;�n)��5(?�ۈ�����p/I�+�!L.#N���#��G����fDn;5}o���Z�f�-6x�#�1�����-����7����j���q�xY�z�΢�R��GB2k �=иfZ�h��a�_��7���	��<ܕ�����zqܴ+��ݐ���1~p��̶6��� ՜�}��8�=��-��u��?��u.#�OCjLe#%��( vs�xM�-8����%�՚�V�-wXV�5����W�j�ɼ�-�6���2|-X�N�`��h�� .hXF1GD���J47�^2��s�Ě�EF���XF�9�U�f��.�]L݁˂n���"& ,#10�JL'��A���F�'�(��Ja�BY{�f�_��}��w�x���E}��y ��m��ZJ��!R�]W��Ww�>k���h݂�l׃	M5qH��-AD��
d����D́��=���n��O]Ѷ�E�kʉ�W�|�J(z/t�b�)�k��D2���P\e~1��#iA��*7.F���ݐ/�Ĺ��,"G��Du;w���Y�X�4��-�@O|��Y� ��E�邖�Mr;'��g�L��ֹ �.�k@�720����"��d���dՑ[�@*SG�C�}]�Iw1l���M��e�@�%�`�Ѩ�^ǝ�nH&b?u#��P���F��{��o����-@�n2�[R��Y��9ba��PU,F ��^���T�赠�ĩ�͟�\}Tmg���C���q�_��(����~��f��&�t�u�9�BB	󁹰T�i"n#ua�P�|���&>�,��JD��^��l�ʴ%=WjM��R7�v+M�����v ՜�Ӭ���g������]+��U�d�	9�a)[a�p��+��bD�K�9Ⱥ�_�w4�7[��I-��"�1���1tr�i�II	D�/3�-�6�d�t���p��ѓ�tE�N���q��-P��[���hd1�k��i3��B����0)�����8��Y��'�l��	ǣl�2�UPH,K���OU�	j�xq}�����>y]yd��h���S��W?N�?.�5���:���<�$���%��ϫ|�@�݅�X1v�*rrj�K�L�b�Q���j���X������9I�aᳰa}�v�Ib5қ�m��b	W?�#&���?�Q���	2�-oE`�	�K�����N플��������]�e��ʑ�`�^R�$���d����:�S��B��]��I���)���8�aE8�E��ʁ\@d��W��T�D1���=c��뤷�l��KX~���G&;�a������~�(��kbI���^w��T}5�>]�imu�m(CG���圸�\����o
�;�`_Yp�HY�"�Z(ŬN���Yg�����<�.�	������F��4̌tY][����E��3S�8E*�$����V*d���T�������&�n�)�d�Y t�-�@����N4\�=���g��H?(v65���KY���T[69�� 98V��:���TD�����[W���Z�ҊAU(0��f���, c#��BL����
�h̘�{fy�"�Y�V�c�.�:�O"5g��dK�M���fVgߥ����1��\�>r�O�����qd|b�{��B)#�\�.��%_��Xŕ_rcwy,��h���~a��c���Ũ{l⣻��_Ţ��.0� T�?��:�x���W��e�샼��b�gss��p��URb�_f(I+�6�c!cwb�ޡ��()�뼌�%\��a�	i��s݌��h+��S��`�T�0;I_7���ULF��Z������j��i���`�58�Q�����)jۚ[�a>��p/���5?���a
M��6��c�B���q�GĨ=H�N2�P���RE��
�)ĩ���4�T����q�	�H"����´hM��������¥�".�=b}��q�t���+��i�v@����V���
�w��+�A*^�ϼ��O�e�"�%cyo\�/7ϩk(Y����������]*}R��	f�L�Q7Ǝ��C4��8���}���t&s��u�Z��^��Ƿ��UN����.��k\���C�3)s�V��vP�:[F��t}�Z
���/��-4%TB�C���~�'*R�K�F���Y��{a�]�������(���$aZ���ޚ�/P6#��f�\�M">$�!N\cD8��
�5�.��y�sf�B�s%�~��]�4Q]��+���=}���9P3�wJr���f����up���w��ʤ��V�#�%��%�}>(r����u,G���2��+�o���/w%7�=%���ir� �5�C���]���:tlA�n� ��E�R��H����������Щ�,l1���w6M3/v�/�;%`����+�1ƫ&�zqo�1�	ޔ����VYO�
��C��?��I�~��=��c�0�&��^��[��h~L/�6z@��@y���������N�]+
�x<t���S�]3>��r�η���]!/��{U�u]�����n����y`��en���JS��|)J�%�F�@��ss���q�,��(���bvstpi�w��4�h���e���Hd,��8l��y�.��p�o|?4	����'��>o�����r��Y��� 1
�[U���-�8zQwF��s,���\OVE��4��,�zhҚlZ�/������A��������ؚ8�V��v6i$��%|?M�V�x6[��D����wS(�{�l�c��%��(�QGK�ěC�
��>�"o�D� &ֈu�b˙�st��5T�F1�d:����N�Y�`��l����A�����S8lz���i�Yf}�+�=���\-_�d8�U�>��](U�� {��t�<�tm�L�S�8���T0�)b>�8�z(�w�G�@<r�9�j[������Q����`�N��f�Pa��WΆ8�Elς��wW��$�e�՗D��R���v#"<��v'[d�wE����E�֚�h�*A+�uR�&�[9j�u\1�(����a0�X,M|�.�e��lF7�t?�����o���Ƥ�c0s��#R��i�{�=��xP��㥚� �'�0���{����������ܽ�,7e��t4'õ
-x�`�H� (b���+��Y__cB��6ǅz\��>_K�g;��e�����J���mK7����<<�\��Z7u�p�l�C���d��y#��	�����9[ƻ�G�O�K��©�aD+
�W���$m^�>p@�_�9\�p��ί�:j���ۨҸQp��������9�zՠ�E�hnpm9a��~��B�Č��fY,K���:�y&�b��m��S�Cn�^e��k�'-����LE|�����ޯ�=���/-ne������$Z������3�R�mA�D#?v ��?8N(=����눙�$�sM}\iC�W'��D�J@�Ƣ}�	!�Vz��d*�a��.��9��4,�)�^
l#�e*�4y�S
3�Y�/���0��`��D���/��Q?ns���Et����䋣ҭ�>�nf�*��"� �2��<�ղ�D��b�,2�&r4�}���������b�g��O@�*�Q�Pe䣱p�T����q:�}*�����!��P&����PH��_�⵮�����P& k������:���XƐ3�愄�&%�'8���y#�J\*w&{/�3n\u<i��MP� �ˤ�R̈́M�P�2����)�xW�����_�}o�rz�g��d�0n¢hO�)҅�%d�3���fzrb(	(�v	�v�f\�D`l!D��bz��j�?5�Ƙн�����`�?��ؤ:#*��0��3<�pe��naTC�sWu��i���IvR�8˪���H�*qI1�f���5�v�~G��iIL�j�q9���K���P��"����]�b0ޡ����'ln˫W�U�Yǧ��oEM�j�y���d�<�%�F�T1�_�v��̷c���}��r�ڠ1�A�Ӆ¼�,�4-ş^��Z:�)=������1�F'�*�3n�._�y�-hYZӾ�&�?����a]�_tl���yG��Dk]M����Aq���_�J_�+�q(�:�p���͛&d�!(}�Ϳ�)c�<��L=�����W�����{	!	���]T�d�4_v,�d��.d!�.�,�mb�rB����:�o��օaC�G��\�J���c��ۦ�q}
��9Z��,���>�2���L�mϊg��MlG(��q�K��m�J�*gK���7�������+^g�"�X ���L��~ޑ�΃t\IC��A�k�Ct��T�5�OM#�]e�d���;w'��mŶ����b,Dr����Ũ%б��{@�'3
L@��s<���fӋ�u��קm�R��X����^���8���D��A����S����X��A�Յ`c�>ڈ�&��5"��k�)��Z@�U_���n�3�Y�?��8�����0k� ����U솾]�[���t{��������O�
,�;�V�Γ��)�L�Qg�9cZe�W�ϲmw*j��6
�g���N��æ@���O��6:EU0k����*�Vh.C�f� �����k\���	���/��ͼ�DJWK�dr���6,W-é�_�'j�"���@T���*��:��~L�m\�S�j��J�ڠ�a�&�FK��M6���|��y���,���#B/�b���/>�w��ϝ�0M3*�a��I����э�(Zi{��f���B/%�t=3F�z!t���
�d��~�-|$;'��s�~R��������6Q�_�F6`�F��_� ś��=3��(=2�����~���{��V�j+A�c����R��Z�����5' ��8�J����������Xo�_+�
�G�iK��Hx�8w��'��:���r�5���>bذ[D�]ɏ�� j�B���Ҥ���dx~��=`L8����zO��� �f|���#mӝ�mb�a����Ϸ1�T�y�}�!��Y_�Vl�v�F}o��c;U��.��k:R!�i�[<������	�D&]�����b��D��JZ�b�y�Q�p�2�/)X}[��h��P�R�����"`��7�8A��������J��۱��� ������Q�p�ug���o"��(Y����%8�b�qo�(Xo�������c�����)���&��FX����A�ƣ��a�N�b�;�P��)�pf���L�v� p���7}���|�`xa�W~��92�W<	�j�u�G�_N�b�
��D��<��{��� ՀC2�GL�P�򼚋�3xa��;�zuD�w��;c��e�d�a/��i��VNezb���2�V����,����������M"�%<�O�[��Q0_Dϫ�X�}�N���R2yg5�|� ���h�jO��2�D"�u��kd��	&����C�vi��[�����3m<a���Q����/��w�8�1�G�@{�x�tӟYl�?"WP����e�FC���7�pi�s+��X����s�l@��P��y��Y������;0[���K'�
L7��`�x3Ӎ�.��3�������p�(#���wi�Z�v��`�,i�I@�c��d�ʅ��HX[r|�|�^OO?wѬ�����vP��/���/�_
u�G���\�x&I�����k�"�֚�2�f�f-΂#�pr�[��ӱ����:�1�������8� ��r�Յ.��]}������p-��T	�l���*�9�\���D����E�]X:}V�k����ۡ՜��}ٹ"��Ƭ	����ě�t[Y*d���8o��sGw�Fx�E�A�󄡺(!�2��,���+V���X��;^ް���ʅl�'@w��~��o�wTgR�!�>㜣������5/�3u&s;���aoٓ�3D��K*c�;dӷ^B��?
���Ot��|��LѰ�\}���">eз2#�龕��֒����ݲP�5�����:c�>3�q�������2��o���$�,�2�W��#��t�h���:b� �7�ڰ[�&p6ߖ��)<��%�$��������օ�r�qM�Px1��� �:����IQ�K$٦�;g^kki�<H?Y��0�1���P�*K|1^�MlS��yS~H�۳[��V�`�j�K-��(��P�S���D�yr�\�f��ވN�gLX�S8=c���1j���p]���'�w
j8}`O^&�q�I���]6���G�ꟕx��B@ls��[��-D�x�y��=��CH�H�%���`z��|����-,юϑ��l�_v�>7�r&��7u��>�#^&�`��-�VE��y`Y>��?#iǥ��>0�:P ��J����DT��+Q/$^�[E	�A�p�q�W�Ї��o:�oQ�p<�; 
��P����Te�����7�Oj�i�x	\x�����i�lɁ8.�����V2�V���
kVp~)�#�(�nC��d��}�O�	w����d��)�s�4b�gl�?ϫ{a��9�s?d��`�7�xf���F���^��������t9c��%,�o�������?�=�O�Azo �F�E4�1�ęs�p��Y|�E�͓����.mW-��f�t3|I�1�E�9�� ��8���$`I����t�R�|��\���Lg�"��V L�W����X}�/�/gʗ��㳠���1���k����O%̣J�ff�"&�D�*��)s��C9�&������m�o�b�􋧱���o�>Q����:5Pl�X9_�ʙ�����G4JVG��{�"P%b�L��'?��fjYEԳ߷��i�����׳���۴ѧ����I��v���q]�14��om��7K��6^y�`�`�o z��41�k7ux���PV������q��O<��I����t���VbR�Սz������7clW"��"���x�{�3ߝc����<y�O��[V��F�Hx�ֈ�	�p��F���$�q8�=ϼpކ�l48CiEw��B"<��m��M%fz�zc��/F�� ��G�N�5��0a��Ow!$���5R*F��d�*���gC��,W8�W*u�pƹpP'>���U�Vh|O[�9Jp��(��Z�������:���=���
���Ҝ_l&���g� U�2��`3o�Y�c�4�u�OQ lrbm��`-p�y��}�=���,���zZUQ��:j`l+������B	�*�_��D�Gև�X��Y�@>��*D�e�A�}�(Ԧ�����=�W�2�t�>�3���5��C��HN�}һ1��% ��Tm@��O	6��
�������zAn� ���O��xi�-m(�"��Rzl8�c�,�$�+�j%����H��t�+��#u�<�$�p��`�	%?�k%�	2����A�T��y��������U���fC߂�xy$o�;�R.�GŘ_�-�>ŗ�S 2�x9ig�B1�bǪ|��IT�坩�qI4�$سM�aƛ�'&X���q��E��3v��l��wC[3m��)u�ǜml��N<na�8Nw뵀O|잗�ZKW��'$���I��	��A";Q3X���5��򞣩��K�c�\�Ѕ1·X��~pAM,ss��h�4������Du��w��'g*T�j�	�'�����$� �֎"�Q��T*��>�3�1�������y�4������棽�ί�������Iɟ�Ʃ�ɝ�b��h�����'��S'�%�ԔD�de�O�xܔ�&���r8�8��AS"˛�-���o���h=8�ci��\7�\dDCћ{f��E���#���m�W|u���^y�H3�I��<�G�i��a�;�Ù���@ؔu���@���֢��_�7�7g�W��[�=,U��8��	�e$}��)���}9_Qž�.���mV&`k�l�qT�ծ��$fE��}��\�R�Ou���Τ\ꀷ-���U�}.�����ʟ�D�&F���]��9n��	H��&��:O��.]F���x!D�τ�Ĝ(�1��<[�n]N����dM׳�%��e�a�6%g q�"v�>����`�P���(�A�^����<-����7���5��8��hc}�?m)�p���!}�N'=�T��
�c�Pl ��n�Ժ];W�����.�9�&p�u��2�"Ρ5c>U���<���Bz@6!u%WE���m�W4��x��1>e�P��&��k)��y������Qlÿ0YB�T��>h���sZK��c�-�^���KS$�d� a�sd:��l�Tn�m���U�u�)J���F͊fWv�X����K�I��H�Bg?�!qȃ �i��9K�W�A6�,=����;QO�ǫBq�u����g!7�P��k?�0a��7h�іW4t����O�?��m��,���t��7������D^}=`4N_X�������u9�@�<�}�Y�ZsAFɲ��1|(/B�/�ml��1ɒqЫ�w�Ǟ��9��rۿ�q��L:����^�� ���70ꐾ�36,�w�9��S�xUK���H�┈�s��gn��N#i�n����� �i�����˝x-�9�A{(d1�<0!oU�#��CVSf����S�}ju��K�k���qR�>�Y� ����E
Mf�e�m��Vɓ>���R����I�B�$�8w�*�]�ղY2��|'��,x��q���9���0.�a|l�����j�0h솧I]RN�N��Ѡ��Jѷ�x������=]��qQ0.��_o��=îZ��D��W�����1y�|'�󺗼e۳���.�fu�ܧ�&��y��|G��r����c��'�a���x�p�{�K_q.���ZvY��MY�"�9�&��ږ��@��PП��- �5�4�K��&������g������Y.klO��Sg17�6�n 3X����8� 0�$�vZ���R[������"QJ n�&�AO������ƴ�0-G��Z�n��Xi�����#<�GCJ��hwM�Et�-�h���,kϷ&���Ll�F�8Cs�&���L�e�����V{�{5[��v�y��,1�
T�����~;o3ݸ�`U$�ݴ2�ɕxpPkWy-�gYwe10�߫DR��T�M<TI��6ujQ�7�9�����,9��=<���:�j��#���X`-�tnl��n*�vG���K:Aqc�8�����|D?�X�y�����,���(ׇ��E�
�d�J�����iIa��8lGi�����E�����)�ѡƋsC oR�,�R��?\R�iڞ���ÿ��L�ш�����9�Zc����EF�b��@h~���i�:mxR��>�/t���X�TG1�Gp}G��p W�\К��!$¿��1Vv��>�����RT@(M7��̛Vߨ0̦�,�Ig+���\G^��r�p^H�;��g\�l�k_��<��2{��Y�l��� 7���}��ʩ��Z~k��|�b��'������9�x��z��	���nCQ�C~�U%�w�N(�l%�:�s�P��T�	k���	��=�c�\��ڈ�-$)��lV��[��Rcz���ma,�=�]�Vr.pܯo�+8�$r�qYۿ&\����ܴ!���9r����f3�����bЛO��M�{!eG���+�.o<3
Jŵ�ܡnpH�y��DG���//go�^�Ao��r\N�*�4+у�х̙�e�A	+x~�ŧn�%�?��W�KT>�$jq� 99N�׸�`���m~�$�仧�Δ嶱�5[-�HR-��)�|��0�v
Y��+��_��)�?�/I��ӯ��M�nE^��k�6ij=)ꀁ����Z�h���w~�Х�T�'���;ޚ�f���KA�/W^vp� |������/|�Dn9QI2�=�X��Ӵ���|AC\md����i��^Vcy>Mࣇ������}���(&��t�la�����+��@��Z��N&��]l�/�A8Mɖe�7���/ZYay��^��!ޫD�0uO����p�EA)���,{n�1jO��}ܿȧ���yPk��UtI-K6�~�Ժ<��P��=ԏ:p:2�4p�!��H҅�M6� 0]v�N���F+~J�5��*�\j�T�_�@�}Ƶ�6�_����6�����)���ȯYjC�_�og��Tq����#0����؆_�u5�$�)San ��H
��z��}|)�AO0Wv!m�=������䯝}e����3������^�U��魵"��uՙ� 0�4
?���2�J9�	n��mnr�Fb/�
�o�!��44nLN���4�}#@X<���à�����d'���W��Ef�({�os1A^T)�c� �(��&V�E��!��L���a����銱+�3�#˦:���ѷ�K׷-�\�^�L�>�8R����fl��ĉQ5]�0lOù��T�ý�<�!I�#nUI�R�_ש�~�}��q�w�kV�uP�}-�Q �l7���딝�s��}"9�����ӽ�ì)��@r(��O�?P+*���y�X����Q	��>ҬG{̞��F
a�
۽�<��B���uh��� A�$5���r@�#Q�ۙ�6�8W�I�+!/d�Q)j�M�u�yU��?���5X6�����3��+v��_`�aȀ��>��	V�#�t��P!��R]�l��mט�:�Y@ؚS�5Ok>��N��!c{Ğ���X��/�Pq+��x��U�"�6(�'���$1�*z����ިuF�;5ؔ��������0h8p�;�J��0���N^�	v�ׄ�_�Ô�C�=Z.�>#�3,�uZ�K�X4аS�������qhك��=L[�q�t��Q����\���0곤O�I�t4���NPg����:uc�� ڔ+��o��Tk�u��0�����6�����ÕIF�,����l��F����սtHs��wK�h�-�+e��=�"����S�a}d��Ś^t�I�Ӯ���m0l��7��L.�TѮ;�u�|.qFnc7Is�0K�s:�?�I�53hPUe� ��➩V��sJ��ί���2�a[}-8�G�9�� �J�G�I2�81���?rt0�r�nnVYcF���\%�`����X���Iq4�!�TTj�$����0���)J[��J՝P�n:�Y���Oȸ�sA����s��'>�h�1�fG]گ.Sq�C�B��%�2F��J����Ь9ۯ�ۭ����"Uf�)&�s�u�M�l�?�A�����r���P��G�K���S�\� ���$��N"��2�〛�����x�܄�i���@u���+���=�����wI Z0�s��Z����W� ײ�B'�`:�=Y���Y��n팘o+sa@���"��o�k�]��H�j���S5$��2a�S7���#�L�H`S/�W�]�c�.����`�#�^Ij:#'~!�$.	oê��8Z h���-"�Y��gKMGei0���T���x#��~�K?:I+_u}��K����[�a��<Y�jZ/�b��J�u7q���V�#͝џ�x��,�S)�f"�j�=}��P��9D
�	�������ϲ������L=Bo�*W�ń�2ĺ/�4�,`�n!,�C���0����ݢ���-���l��[R�^&���T��f<�ۙ�M�)�=�.SwqZ�or� !���)��ה�����ߪ��6_�)v�%������j556��!^}n7Q�!��j���Ji�l�>�0�?Q�EY�Mm��kV|���?���]?�}�OUs�n���K�R��9�+� /�7��%W��\	Tչ�``nԈ`�>q�'����B���YoFg�H�"�q4���o�G�����p�w����~c]�>  [ƛ���CLᢀ���Qg�s҈���x����ew�d����ф��;��Q�oo�x]?)3豃@���[q��	���^;�K
��,�Hl{9R9w�7� �����
�4�*(�Ca��a��pya���wZ}�l���ģ��G��K���ǝ�`!�4�"4
bfV���u,mAp��(��$��q�	��D'�9Z<z��H�8%���e��QZ�w��i������&����'�!�NP3r������k�b��Fj����arW9�}��o�N�E�����/ǖñƾ��t�6����ɳJ��fY�MW���%\!i�D��֭��^�@����3�����|�C��`�ح�2C�
�~k݋��E{E���R��'�s+9*�Գf����,�f�%}+3z�V˻�t�2L���NZ���E�l����dC6z�B���Hh=���Ȧ&����A��4�E�z�aF��k^'A����ke��=�7
�]!���������π�.��«����"{��k����P|(a��,�Y$SZ�O�n9���D8�<�y��d*�{T��n�m���3ϖ��ί�w��4/g��@T=��x�?�[x]�<哷J��-�(di5���@3<�?f���Z%���)��Q�2�HRp��V������Ӛ:B�	C� ŏa�t�U"�X�}|�Ϫ&������o{�+��ᤰ�G�	:f,����<��v�� Yp���ձ�q���̉5��l`'����wV͸ê pMc~���Z��-��nI�����W,T��N0������ w��P�)�F��?� ��{�T"9�Y���C
C�J�:��Hÿ���]�)�{�X�3Q�$<����B6�{*�'���H�1	�����/�R�ܐA��������C��0H����a���[��Vo���Zg�f� g{��/O�o�2�3r����_&��I��΂�.6��t����4�2`��=S���i�_6��k(�Edճ�.��~�q�����F~rnO�m�MTG$x[�������B�j���z�������4�D���b�J
:FR^�(o� ���=h�$�� �@�H��nx���	���n�V���b6滓��д�G�rR��-�[ǽ��m|��m�����m(y�W����6DLUR��4�X����\�1�·�k��T� �$R�m�)Ug���^9�����;�[��C����5�z�C3�Wd�Y7��-��옫�0&�`ɡ+���8�(!�$J�)ߢ��GR��~]��B�m����J�%C���D���E�P2DvY�ƳOt"��<m�(��#��7JX��]���h����9�Z"��o�{rPaQqn�a��'ڪ���Gү�U`z�-��>Vy����a�5�4$ڊ��FRմڴ��kM�j�7��u�mf ��)���
�t����FЮؙ������xr���Cׯ;��)�<RS�V-'#��h�e�G�|y��J�=�U)�6]������x�v�|#��|�j�ɄA��P���%½�^N�2,�W�/gH�� Z�������
N*���=`����ɵ3��+�a�kJ���t-���_�y��4y�p�m��b�K�j��U;4}�X}�H���[� �,�n�ܚY8�t�)a�E���m,�E�[,��4RaH�Ϗ�i�����t��?i�}�\�`�]O7���Z�/*�yPO�)�x��y��Ka&����������!Q҄��>� ڪ\�3�p��ϣ��Ae'��N�Sњ�iFQ���%Y����
_�}�2y�GV]��cە�=��������HB(���#�E��~��S/7K��N%�l���X4g�����ċ��3Q�#+��ڇa1|�`����{�>Ļ��x�3kׅҩ�� R����9 K��PJ�tF�+������}<�����!P��PݢÄ���q57Vӱh�Mo� O�d02Ή�#G�j���C��	���Z4J�ҷ��`�ϯ���Fv0��s	�d�|R�!9��������:���īi�������l��S!As��1ǐ��UR6J������c�
���Qn�8i��|T�����ؗ��qa�`9VcaZ��P�)���P:�V�lF�
�����wQ����c{�ۛ_-��e���G�!��gݬ`���J�*=!���G����Ai�ĝfx�-��+8���i�P�nw�q���5�S� !�y8О�e��]�kR�/Qq
>a��,���l�cPA��>.��p�a�kg5G�r��a?Q�&aS�ɂ[pB�iSD`ܻ�M�C�y�pLy�,��g"��g��%��$�@�o4�@mY���u8��J�@	�&od~	rT����[�����Y�.���~�0�p�շ:A��$`���9�߾^�*-G��O�����Q����$H�jGt�,��!�)Z�F~��rA�W�W93(���w"ԅ�9�ԇ)��s�!�1=D9 ����v陟0�8�2꾼sQ�Z�k@�J�3_W2�1F���ю�'kR�Z�pX9Q=H�D�g�������dʆd㜛UC�E�3��hH�G���9�;��FR�6�����넝���uQ��!�s26��'�}�N��*�}Jl�Me�u�Q�������P������w�J1p s��HF�*����L�$�U�@;���%?��4v����OF����ͩ���_�"��x��;�64���&�|6H�`���%[z���^AY��)�'�fI+nJC���?7�鄵����ʑ��&ݎQ��W`@��o�U�kBo��9K����c�:��T���|�f�P��X�h
 ���&��7�.����N>�+�FFt*�_
���Ҡ1�{�h*�-oJ��R	̲2���ʍvC�M�R�Ƈ�,��MN����n�����g���Bj�o@�X��#+��g��e�iO�F������HS�<N�qH{�Z�x�1/�R!=o�(����6FÐ;��y Os?�ۑP_`I��|��IB�ú�-�J�����||Qo���D~T��xz���t.�����Q�%��a�2��DR��߰ ��{����f��m =gOd4p���e�#�hl�=S�~�� ���������O�����z��J���]֓��b׼-����������{�P�A,���OY�ܮ����3je�Z�){3�q�=�7�!��{�Sj�\M#;��v5E�*Ug�i���+!h���٦@,���[�E=�O���;�c���˯�8�.]6�`"�q�ᆒ>.��%�۠���6Z�bЌq��v����R�@�,^茣�ԫτ���h6^M�˗�vA7�����z5<�(��a�jL͊>)+�DV����>��1���r���
�8v��˷{��=�������bF�lN�6c�:���=L}_�[����47!���}J���/<�R� U��t��n8a��G�NZ�S�M��K�~/�[O9��*L$Y��p�J�O�Tŉ$�F�ڠ~�
��kΒ��%�B��_�%
<�[A5|t'�����YC�0�Ǐ�.�nX��v�،�pr:����ͷ�����[�d��Di�9�YW+�H �4���b�;��}J��&�de5�C.@�0L�	[��83:0C©٦2U;W��;���l��� �����e����'��r�-l|sV�?w/�^ä��I����<(��C����0�Y�f/����/&C��X�^n��2�F����.��%-�X	�i7	q��6��N�}9%�R\o��T���`\	�q��%&$��߂�4�`Ӏ�SkW�ɍ
jVD��M�#���ƭN�X�&����K�~�0�0�<G�v�z���JVp΢�E?���*.Ʉ�P�&����2�\��x�YB���"��W�o�GNQ�-6;�G9��.�,���ȳ������y*��I�m8+X|Fj�6b|���wJ����H�:���9H`�\B��.G��z(�����G�#F�U��a,����!��i�����"�v'��^��Q�%^E;ix��6��2�S$���_)n��7R�(L}�?�(�f[=:YW�������ݴ-�]����1��S������'�<e��XQ���ej_�b#L�/�-6aP���m�6B^��;U
'��J��1�+�q܇8����{Z�LiG�)���櫷[)�+4*�D+*^����� /*�G��EƗU	R�kA����>�܍�A�/������.�١��-��W��ϸf"��/�s��������v�Rpx{,�FY����"�UK=}�79<qƆM���HD����vr>��� ��)&�M;��GU�s�t7�s��q�a��t&I[X>�kѥ�� ��@|kĦ�T�\0����������yw��/5���v�G��fC�	���<*IǞ�u����+��Bʮ~s1�y��;F%�g�Q�r��$J�F;ٸ��kю�(�N�خ�m񆴱��RF��^�mf�`�A��+{� ��;s*	2&#����!�Z��:��ߘ��G�f ���:�R�eJ��J��1�Ѐ@�N���nb��g`��Ôʫ-�Y��������Ir*��K���R0�9�jlb	�L��Ӎ�qu��W�\n���o����v����"8�*��cô�a�(vt�
0?��K��nI���A�چ��=��(G���O�����ɹ�^Ug�[.�jJ��{S��"��Z����Z�ԉ�n�����V�1��l��Cu�Fs?�=RR'�1������ǜl;Um�3��L �-��y���gw�����7T�: �/2��0"������]�Yg�~*�A�=���U����$�D�W�=/ ����M��p�0�;��.R�۝����@���F��f*���'�un�O7��4�/2�-Y�#���}� �D�SZ��X�B��0�3/
dq��MBt#�ۙ�`OO	�W0Y�;H�ޭ��P���\c/y�v?����^��F�m��������g����Xk�"�u5��Z�ل�<tQGE"pz(��e�&�qq��K4���}���x����B �b6(�� y��r�_++3�(�Gf�r��I���{�襧*Ⱦ ���
K�E�8�ǵZϚ�rs�����*�
��%#r%iܜ�@�S�E��>��b^�㪅�]��e$r�1���3KT$:����)�q�e։���ӌ�h4-B6�f����b P
��	x�:2*jxɜ�����3E'�o��0%��C8]ԲK8���߷�i�(o�ⱬ�e�U�p�@5�e&�����*�6��\��%^qm�7�1��������)������-9��0p�u�N��SB��r��jxP�u�;��:�B�|ގ��\�������X�"�t>bO|�"��Sj�Y��6�f���7l����p�������N��l�[0N���r�f�65�*_4����גMc"��ܝ j1��n䠨3Y�G�A,�+9ԛ��@��9ݴԸ&{N���z�~��p3��������?�+���Nvu��������WpZ=����F�m�a]��5�ѱS�O��mE��ʡEV��8�Ǯv: *��x�F�s��~��S�k���6{IU�|���kv(D���+9��
��nB��E�����lN�=J�������ڂ#>Y܁�@4y7"��$���O\:�&�՟'�!�
c���c� �$x�IHz�U#./��;�k������U�*Ӱ����8��A#R]>�i+�dBs�.�{�5\��'���؆��J��#~)���j:og�5�k�&R�!n��İwq�G���4J��`!��O�qc\�d�/17�K��p�$�5-M���<�����u���&G����hΖrجH΅.0�**�O{"�l+��k+�NY�>������oR���`Ҭb��u5[�N=���R�B��_n)]��?c�5��Y	����&�v�>��v�
d���*���+����$c�2����JX����@����Gu&���atm�s��:zY-)r���䄯��Ͼ��5�n�ǈ�Y1�E�TӦ(L�w��!G0Γ��ݣjxp85>�lm�%��6��
�3����~�Df�ۖ"]���Oq�$���a_��e�(�<5�[�+J��3�X�����ҙ��u�u�ĵ�T��1�B�c���m�����=�s��N�u@��;$�Ni5"�	y:���<�m����#6" ��m���$^�/	���r�o�S�G�4^jz6F�*����jq��M�2��"���'��9l@�4��~��{�pe� `��a��C�5��VNp£S�PX���*5�g[�wa}�c��^F)�Y'�j�5�)��F��S#�u��mw�v0)�����U�V���&����.>��Sa�p�%,Eb*��P��HC�]k\yq���@�41�2��Fw5�;9Q��v!�J!VF��T�C��3#S*�^�,����z�0�*��.�JE�3��v����j*��*1;�6.�A73Jael~�K:���{�`��h�l��R�:�7��޳D�Q�=dj�'{Cp^a���DX�^���}F|��t�2�(�����Sp���^&��q=��d�t;�^�s�� _���I��G���6� �5@�V>+1��i����ċo�{�=�E���=��,d|k�i.F]�RY���/�����?�'b�yga�>���pem~�lh2Mbe��B����X���^NJL��vm_djb8|�.o���j��]��E�lǂ�	Ή��43H>z1w������x�f+����Խnu���~�-rU1a)��OnI�?�e����P�8p��L�w
`�.�*�����@���uD��;O��Z])��
����Ys�����@���wHΕ_tI��aNհ 3?��:�_��F��pE놫ʌWM�?p?���QV��H,,�i/�r�e���Fs̳x�a8���\�w'��YEJ�&s�CPt��A�r_S쾙T�^re�s@B/R+@��c���)î0�,*��jN��Rni�@Y���iT!�V5p���ϔ�����Ia"q(pui*������.��(-��>r�y��{�N_�>f�x^��0�jҰ�o�����s�Mq�#:<dj�x#8�
Җk���%Hc�k"��Cv�,��`�P��{cH���@�&�3�l?�-����Y*rS�e���Dh$�fI��X�D��

���̟gݷ�B��ܸT��a.�gק=����2ȓ�����L��(�T�6��>��,��8����U�edv��ݚ!�o�oϧ��)M��V�o]1�[��CX�..>���=c%!h������3��p�+����l+T�:�뷿�[�k���%��n�O5�F�U����S!VTL��2� �o����	LE�����b�a�p��<�>ㅏ�)�V�`�!��d�����#����X�$�b r��yqwl?�����0.�V�#�Sǟf�tݬ��_��G�e��������!��&M�IU��Rk�ЎW�ʴT�~�� }�ep�gTi��B
��&~͵���h��SW3�@j�V	�F�UVU`Z{ ,�?�}�QGCLR8t-M�`}�J ݛH%�(Mzh��Pދ!8K}�5�(��� ca�4��>��yP��P��J��ם�2�"�73CH��<dF6r�0d��؝���VLQq�v��v��;n���������q�t���\����)GP?�˻��%��m��0�|�_�H�'�JwŶ��^�<�<5�E�H?��Q�l֋ˉ1M�:26��&�F\�1�yo�H~>j�y�-�@�<�
��O%�]�H$ ��O�w�v�}m��M�h�*����z⩤`�ʌ᳥	y�N��f/�����y����;���1I)�N��~����]T>�9����h�<����\�(o{�#s�3%r͌�}l�Z��:���g�3�k�O`���k�;��k�bD^�n��A�m�}9qaT�
���(��)�G�����SR�aX���2E��������,���aEO0��s	���O&B�P�.������k�}ѯ�#�5@^���<�sn
:v�7UA��W-��u!7�M�ǟ{�C�2UΘ�,m�;r�;�(�fa�gF�^?ᬟ����0�;[��ˏ4V�"Ll�6�}��2�4�iD[�{M��Fƚ��D�^z�o+����Z=/`��t}`������}�ʎ��.d�0{}7x����f�*s��~y5>�`��G�;J GH��� ����P��﷯��lGȀ���+����j��o����WV}��	����c>	Q�#�%O�ki{KB!��}@S(��Y����wI
ˈ㩜�t�ü���Pa��L�~:$���$_
�ߝ-"� �	��[��+� ѣ�T�HZ�r�9_"g+��+γ6�m==�����	}ٝ�}�N�b���s���,�G�Me�!�%X@Ƚo�c����OQ�tߣ|d.|C��g�]�xN}|��_���0�������Ɩ��4�u��M#\��`�9#gR�b3TRB4�^%s����~�W�Q�{�#)���J��v.z����)ӪG���f�fkB����K*���L�y��z�%)�:�VQǀcV���Ggx�g�)#�]��e<㍟U��[И���e���:�6�����Ʌ�����3y������eC�¿�� ���2��xۘ�Y�D��R���~&�2�VKͩ̈́�0�#�ې�<�����f���N�]z�Wk�T���i�x��v�T��^זۑ	��Yd�-�+�����g�dU0���RY�}�����C� ������-𬏑}f��"��h�C�Z�b��v��2��lG����+�w!��j�JC#Zvpʎ�qr�����������9GMJQ��/ �V�>8�CܔW�������
��CYrlm)7o�LJ|�-�Zٿ���<+�ҥ}�ql��Y����[-�;�2��qo�k�l�[,���M�1�;��?�[3�^��h6�p�2<8%��T�,��/޷޶>�]�_�'"��&	��������OH���>G�'�<�i�
@Q&��ͽ�x7��h���������~c�߄�.h���L�1��~L����_шki�����d�ʯ�k|$V$@3�����M|MQ@o���R��D(�`��T�Ӊ�5%���E�`]�Y�T��o����K䗢�� �'+͑Q��Z���l��m9��:Bf+���֐j����N���[Yvq[�p��#����J�-bm���J������"{ ��h���4Iɡ��p���nt=\�����?�G�l��U����>I�O�i���D2�l�o�P��W�|����qS���-�7?P�>q��{�{��6�����Mc@2s�6�-��ԎmF4���q�H��Q�ۼ*�_�}��딈�*wM���&9�H,��K&w7����
46���yH;iK���ݺ��#��A�wD�����бg����A�JvL����#E��S"UDM2�L�eez��B�V�fL�^+j������d���+�d��a�lT��M���7�Ĳ!��ӏ�!�_��(:�b��V~����q����/�1��?��vG���(�o�(�(s�ȕ$�ґ q�Pl	Q8�Z���4ip-?��~D{����,"-01R)��T�RI&�'�^���nM�j.�+�;�͟� B��^6�
G�~K�Ó	��7��Niy�}7��Oc��V*��4GH�G�<��qI�y�Ĭ�d���\�R�[Ŭd�&�F2%n�����vCp����"���xDHr��E8�YC[���~-��PjM5-3���VQ߅���2�Ocʚ>����^�O4�P�C1�P�~�L:�Z�e(���zӎ�;��?Nh����_�-���Aw&� ��1�T uC���/���/B*��q���7�����&@��M����v&ި��Q�9z3�pVd4⇖����#r=X��R��B�_��f1G�le�"	9���ʓ�;m��/6�ѵW�#̧���o;�p�g.Q��=�!�!ʪ��ӻ���RS���ȟ2�A�-e�ލ3�(%�όb����#k^�T�$4]��������>�X�]ʞ��w֞���"Q��\�f��&��FWȆS���x��L�T4�a|����7�D���-���z���0�����ђ�"�`��)��gI@�T��C)��e,�	kp�c���NI�np�U.b&]z	�Z�i��
�@M�]�"��{6����m��g�MJ���a��>�H�se�:������ R�g��ઌ��{55�!
n���-����|��8sj�x�70�Ȥ��
�!���I�[�r��:4���&� Z���6��v��S�[�F��۵��D.����]Tf�Qo�g��]ܦ P�$�Ӫ>A�� 8��s�9Լ̔�hIBf�9v�>LQG~���	���XNiC���:���ޥb������{�hD~���_�ܯr:��lbPۇX�E��C���A�ǰ0�"#`[(ob��ϔs��ǎ�x�4?�/g����;g%���[���Z�-�q��F���hf�{�bh�8{����0�5�V���U-��㧩�0�g�����?1$��R�n3��
�B�B�23wA���\�[�ߡt������|��ɮd�w����K�Tq!�6���R�\'�X�m���B}�6��ĨW`��qw�+3�K��,_�UsX��/4��+z6��}����Zo����e�"��q\�v�պ7���a��R�S��%6��(�DE������S����n�Yctk���[��	����U��[�iq!E*�j�P����a7�u�\@�wO��[��g�f(��N�j�ɥ�U��eB����Su-��w5�\���;��ח��wZ����Ewd 1-W۶H4�-���nJS�-Zz�,�%m��אA�]�8�yc��4� rO��� �N?qN�s��>�Ն�z>�}����;�PN\��KR�e/_yK��z��bV��}��X�9Ɖ$�v�J��q9`|3� z��X��c��(�m�Ǔ�Ջ:^1���/�����C�Z��Lr�w�$����o�C�5��	wʭ�_�7}�D���j~p�8�W-Y �<x�i�,�W��-�dO��:��mu���x�����da&� "+��v��O�,��ȴ[�`>4�e����>��!F���(��?��7�6��[5(ط����遐M�t���oo��=α\�c) �Gr���LpE��w�v����`���׌���ңI��H����tLْ�O!������:χ�_�a�}�p�V���5�\o�^Kn��շ��UN!?g_ɿoʂn[�~�Ѫ�Y���N\]���xj'{_崺�@qH��T����'�Nֽ���W��L�p�5+��3\�5��KͿ�~�-.Ը�
-:��,r�O��T�/���g%x��%|�BZ�M����o]}6�ŖB����xW����w�J���~})d���h8�5�6�rO���D��k����<5���;��|]q]T�"�)�bW0P�1�ڣl�O$E�zC��*ꜩ�Yc�%_�y�Ze����i��\s�f��������/�쐩u��1B0ΪfqƳ�ch�Ĵ��1Hy^�D1����ep;Ed��^�(z�������#Eo=��	{����H�?�;�I���|q�č8��d\�H��D�$��KS�aq&�\�Prt�e�s��N��K�޾:Aw x�w"����TDl(�e]��1;������z���(���,�+����w���Eq�z��Hu=8�����*�@<�M"9�Ja;⳷�m\���eŦ>��t���
��<��T��	
�/d�őj-8��vW��\���
�!�kH�\fk4U~����^y�S��oNB��*v������O�ԡ5��fDs���ˎ��.��a�3���;@��&�0��]�ʠ���Y����H�}]SL���/�y:�5���͚�k܄a6�:�Y�M�c�2��������ń@�ъ�b�U�Y��v��0�<-��|Mj�ڬ�ݼO4�]v�Ǭ^:%Ky�:���P�3f���Z|g��|��P���ꎆ��nu�J`�u6n�3�Nπ�w�C<.6uW^�FIwZ�Yȅy�ڹ\����6�R�K�nmZm]�ڲ˅
�f�qm��B�c��.`�|_��Bw~s��������\`����<�f8ws>8�<$]-��tF��u0S� ��~z5|�����e!�G�m2>��E�r:�B�e���d�����X�ϊb�4��їE�6-G�Q��BN�.��M�ߛY�|����DZ�0��.mj�{����9L�[��Q�&zU Q1�d^���u��I�۰:S�����#�bX�,�>� f�q����̐a�`��G�H���_�c���_������a|�K�N�4��zM�Z{8��n�\y��l>��m�R,����Uʦ�m-�Kn(�ơR�O�.��/�2�=a�R���`�u.��.X�]�f�>q��O�������yP�ʾpؿ�Qam!T5o�g�3�䂌����t���U��Wxί1��w���f�Y]��L�6ק]��On��A��dN�/�"��wk�����H��=�e2��st�+��ѳA!�(&ť@�|`�J�ot���RK�^=�p��z6g҇�j��[J���Շ2�����S��QSA���T��U%���kY�r����^�Q����X*T�*�h|94SA��������j��8~8��EIk"2���1u{�Gz�S�&�W֣ɛoH�)C����YV���3��{��7M�,�2�eY�L�o�?7�6���a�)����}u�;��L�WjY-��V�iϚ�Y�U�ϥ���"�d�w8O��`$��A�z�t�?��6Hf�ܩ��9*�g�B)D��;���q֫�����T�z0ER�b�/[V8`
�Qv�0��D �u
C�紦7n}�uf���[)��]��n��1��0�pHt��=��§�7 .���1�b���"p�?GдѠ����'\kѲ��fK���}�؆:��ضr�G�ջ����w�OߚR(���ԤR�����M+�ǂF�"�,��xhv��qj�������%f�cq���N������%&A��5���O{�^
�o���]֮�����Y1Z��&�	"c��4T�CԩтB�gu���z�w	ˉ�e�cav���������� gRv���B��ƽsb�_e��xJ١6��)/��Y��7�4R^���N�9kR-�uzl�20"���"=5�O�I;$S�#O|;0h)������r>�Ƞ��e#w#�T_-TU���N�M��1-�~wP:�0�Bl�%��M���yF �zՋ(%η�C7`ٳ�C��>�n�7p&�:��ʧ���вT\�Ty�)l�M����gT��⛬E�r��AS
�.q��*M~��R'���K�Ky�za�?��*E�5��ڹ�'ɘ6����9i��m���9"�^o,_F�V�:^�qE�4&R>����7��O;���Bp��CW|9�aH����잯6�#E_J�g�1��I���AO4[{�*3�\�p�x1��}#+� �l�
*�A*
eU���!�"#k��� �_�1�k���0��5��R$k� ݛ�V{a�a3{�Ξ'�	�p��ȇ��R�Z��e׈�5�E� �32�f�<�����Ԑw�/>�k �n���s���:}��{h�*���ϭ�� ri���vsU�o��Q���)wS�CDs�����8���A�q�9���0��"5��y�l�0Sp�+�H�0Qr��l_9&G�E��[R*�ee�F*G-׎h޸���Α�C��3r�A�66�|�u>�ƿi�_�f��g7~$�`�!����p5�!���u���=�K3�����>V[R��-�t�%�V�X��!�~���?��*t�֨�D4�Q �r�W��?�D|�b��5��I��˃Ǽ�.���,�	�J�p� �¹i8+	d��Ёg�T~��C��� �X��ahє�k�
�u������Q�]��`Ac?��䇋�I�z8#^�G�W��#?. 믎Y����*��F�)�_MLb�"1���3�kbi��/!���/�8'g̉�)}��5�V�ɡ�+�-�J�����;�G[6F7"���,q��=`�U6[�O�G�T	�Tl��uĺF��a��Ji�6�9�N:��E�D�z'��C� _�+S�8������<�:��3霸�Mh�.ȉ��6�RQ�#m+��c��w�ֵǶ3�����T D�Œxl��w���ʚ:�ҥ�Ž�}��Vъ'���)���	(�|���Ϩ�<Ex�,�eEyE����U%x�nD��+K��j1�u�J�铒a׆gW5ɦ �VWc�Pm'��4m7 ��mњE�u�Ӻ��q����ц��`7�y��$�O]�6���ދ��`������9_�����Y+��"���>���pT�'�[5��j��A�S��X�ϯ��r3|�G**e�<V<��LǬ��6�;h�7���4�|���w�:�5EG/T��;q�}
����G�-qu�֍�v<R�EA)��(Z#�I|��c@�@&�_U#�K.(lH� ��,��JxWD��
)��4 ��XNT$�Ӽ�F ;�O�4vE�j�&�"��O8��N)�Y5r���`\C�bٍ��S}��f� 0W��݋՗W!S��a3&���,�K��� �\���\�@e��xUw1�H���i@����݄֠��x��jR�vS.E�+�����y�^1"2�5�h�4�e���l���|�^0c(����t�h�x��W?�]�rg�髱�g��F�H*c���ӂ�ې�bm�Zg�T��
1��!K�#3�Ѻ��w�ʴovX k�������g�0�L�^�MR�rV�-�'ȉ ,{��ߞ7�淭�#X2Ac�����S��H����ѰZQ��c�sF����1�W�LhYm�R���G��Ӧ���ꈇ����K��Z���z)/��^A���{>4ۆ��:�)+��׹?��.���o�t	Q����+�V'%�IE��yq��ܓV�^���2��,2p����H��Z:t��5i�ɮ}�ܭ��S: Ȱ���fK�!� ZQ���u�	�z�'-�0�%�0��QA�fw�7��@P�%%��6K�i#�]����H���-=�6+����AZ��W�ES��'F��'��|R��дP/�X���r��G}#��� ;��?�����z���^��TEف�C�ӱ�~7~�go(�=(��ފlo�N���Fj�ت]p2��ʥe�,�?��|^�w�� L8K:?�r����72m�{b��8��様s�r��d6g�̝)��?�E7����ҋE!���4�_�-�{�'�p�L,Mb�O�Oܹ5��0��F�~�?�k�_���M{ �΂]���d;���2 ix~�B ���]��^Z�K����ԁ;qN=����D����ไ6PU%ď��m���!��5�~:p���\z^�����7)m~�~�$(e<yϺVۡt?�/j�>)�D��Q��^9!�9����7�؎��U���u�����v��=�F�O���E�G؈m0C��s�[�BDd���>�o��#��-�|/Q��^WO
@��=����7��m��k����\:��Ee�N6T/�ގ�exB��chW��j����=n3^��Q��y�Gm�����)�Ll��TBq%��?T�+� &	L_�d[Cz�
���Z�6�Eê ]M�~���y%56�@d�"����A�W'���C��eN�&"�m�@IH�_t���9�'�^ð\��9ڤ=��e�H���͊���,{3"�J-�aW҉���p�}.�9�~˚��m�Wu��zʇ����ă������bS�T&�Xv*S���� ��j�2}q�Un)K��̝sj�k�����rgzrA�8��~�R���P� �!̬7�F͞�ELO^�j����I7H�dT�|��?�6ۚ��ڢ[�s�~���"��`��Tp��B�P��T� ��@3/�#(-�Qw$X�wʯG�GE��F$�,�r�(�7o�@y�����V��x�'f����I��z�pnw+��cx{q�I���@�����Bܱ�s
��� yb��4��B�bANHE�*���ʒ|�9W�T��'q�-~r	U�����������q#�* "����A��-�+����J3{��Km*'���|>H��43���x6۟J� � ��H|k�TX��nK�O��]-P-_��c����)y��ur���'o��a�Û郬�DQ/o���^gU�=���.�;!���f�>�����!B��ݠ�jXe��Q��u�<�:uL =Xb����נ��^a<�0�2�'A)��І#�2�E< C�)�&��Q����1���.�ݙ��&�YQ�6(Ԇ�(Y��M++>�i�g�Dk}��tJ����B y���q폄�����
�IƝ�U��#���oe�,�	�S@d��`&�c�ħ#���Di���?��sl���6��<b���4�Ĝ���T�'���!+R0�R����$�����/,�r~j�c�)�3H���m�R���U|˧&i�{�Bb��o�R��.�(`�U��{"ɶ�6�k����U�m�����uF��̍�U�.^����Hm��}�lD�y�783��:7foYA·��8q$��E��ʭ3�����KVm��)�Os�CM��K��=iM��x��{�Y�e1��43?��	�S��`P�>�����'L�+�1-���H����9hq)�����OTm�4�x�=|ᯊ�!� ����g�oو�t�J�&B����VjhR���+��r!lTց}�-���������sq+T��G	� ��h@=ӑR��l��_:|Ġ�pGfv��M��073#���ﰁ�T=�� j�|���s�<�"/BO�(���|�UBS�i*{�E.i?/����MG��) ڮ������9�ގ1�Be�)�I����}B2��ܳ�d�v�9L�D�����Tk5��Z��4���v �x��ii�t���c��_Y�)f؜gKP\P�\��bǰ�aV���Ų[~��Z�&vEY�έ�^�.b�YcX<Kf�B� �%CE�=5]��P���>�/�p����&�HTu�n>#�5���d��� x�B�NnR�����,v��3a����WQka��=3��h��4~�Q%v���(η��p+�df�~B�3{�?�54����������T��a�ZPh��m�*f�sO�0��s�G�^*���@�_�����ޕ&K��M)T��nǃ���,$
s�q7�q����
>�y��g;���d:`9�C���`��dh���P����f�BW���ˎ����"��o�J��+�6� ���x{'`�{k۔i�n��"[��~��$U�9X*��d1�#�>0��d��ɕ\�ݴ��Ay���7�M�W�H3��+A�����p͠qP�B䑇R����9�
2S1fC.R_������#N����o�}7��R�6,��������:4��2��ks�@��-����̥�����+��:F�~���#��Sn��A3EV�f]7�$��d�#13L!汝�	����k�n����޳]X@��u
�n�P����3�w�Ru\�9��ﱐ?0L�Uq騽�f̈k9$��<7���U��d�5��p>7�̓��=>���jV��n�x�;�m�T�����s�)#8���;9�.V�`u�5��C��1V�#�s��F��J�3)�:��V���X�14m�yn�4���p_���cE҃W��$k��V	����߲;�w�@˝	�G�%����6���^KA�����h�K���M�[���Y��L�����RC�(p x���E�_�Js���1��a�P�qvnބ�[�p�jh��7[~�Zk�n����S�~>e�k_�^j���P�\Y�d�9�]���밖,Etu~SZ�θ�(�']z���D`P"M���`�Hw	�"!�JKw�4.ØP<�Z�◊���&�`�ȔO:=�-�����PMAv����w����kb^��{��l�z'�0�.2=P�8��U14k�>!�غ�9����j;�=�҉d�a�a��<�R�a)	.H�~�Q�}xٍf,(����<�|�o��"��B����������]�;���b�:V��R���E ~dއ"e�Y
�r$f�d1�t���i�#23N��jϦ�@�M�*��_�k�"�H�����=j��frJ3F[4t�B�ڔ1���g���t�pyn|��i:������C�tG�(��"����TGԽ�L=c�^�y��ԼV�-�RխI��m��t $]JM?&iL�^b�ЍW��(����"�B�D�H�]a7 /!���'��*��o���.C�#�L/���l���F�J"�I�6���KY��'��&/JR���ܣg,�%zߪNm`;;'�@BC�7��<&m����*5�q-� ;' IEHG�n%�N�a���˪�W�6	b&�B`i���%!�a8��x�<ע��W�RP�G�r�]���U�J}�)�gzx��k[� ��6�<�+���s=�bJ�F�s^=���'�o��'�S�͖�v��v�b&X-.��ܢ8���!���f`xU��IK��
Z�J��o؏�7x����H�;עݡ�N=�ny�G��yKr�Ge�A�ϋesa�܂�O٫���Z���r�2���'�l#Ԇ�$���������C� U��u�A����`���JY+��}�N-^ "{�O�q2FT�4��DS�5� ����/��׆g���OsHl���oЮ��-}I�7�6G~45 ��+�ljP�{ M"ˈц<�lA<�����/�=g�\��3��U#B�?��p
�JLԖҜ8,������.b���}�Zwe`�$-�I�	�8Ɗ�2���dں7΄$��%�r}�cEke}�`F�cL��=̦��e�u`,�z���L"�9u�Uod$�rw��4�_'��Pc�dY���3�`0�V@{�'W�����@4V�/�EH�mL�0JƂ��/�����m	�H�-����YgBv�a$���0 �Xc(m8���yճ���!K�Y,�9]��z�\�B���Oଭ����>F����]�9��F�[�7\�=��[gz�	N�wN�#9	��aXSrt�\��7��bGkS���2���o���FEsZ�d���_KM�,m⡯�gr�
�'9|�ߐ20lU!}�B�L(m�>�y��2�e�����k3�bN/�9��Pߡb6��ʧ࿝�\���s���p�64�1ʏ��;o^����Fg��2��_����e��A1z��^rV��L=�;"����Lf�1{�M2;K�V��l��µ�-iF�ԗ@
�k��Ee�ިf��6�D��5�����qjb��w.M�����nј"m�=����0̃<:�����t�E<�Ȅ�bY$ G09��b�0g?����x4�0�U-/C��@v���u4�)vf.��#��h����L��.D�Z�o	�b$�/)9�܈/֙�-�`��T�@u� ��LQ0�j�Z�F����z*�����Y u�2�eOmEE.����l�����y��c�c��}RiDT{F�t}ϱUn7��3�O�0=���3/��\��R����{�nFr�X���݂;dy:��ͭ�?8�Yx�}�|���孓D�}��<�ٳ���ȠQ�I]��4iv܂�0|��	,�%�,H쬅:֦ VI�%����f�$�_!��A�Ct�����}�26~T�!��k_�D�]��Zd���<��g\r^AJn���B�F"�(���2��/�� M�Q�ل�2=�������+�l����A����7\�=^�te['3�_������2 :��V��Ѥ�����BN�;����Kۜl�WL�
��!��\]?��]�_�y��o4MxW�c�9;J�ug
3(T�KSI��k
Y]��հ��ŏ�Y��3���K�8���h���P�V�.Y;��2�ˎ R�4���^��!���I�����Thу�,��ZOP ���;�3#�� �oW���4Y� �8P��j~������#��p�����(a� >���>�^��g�5����B��1��x訩��
�0Mpl��XOZ�/y�%"�]���{����h
C�=��pμ�K����� �������u�P�|��5�z�w�!͘�����h�}9,B�V�D�A,}���r��~PJ�^� r��=�/�߄�! Q	�#�B�?�;��_���k�^$�R��*G��K+��Lt,�ҹ;iE?jX�d��T^�k�LdܢSx�Ny���eo�NVbvu&�LW���3;�Z?;���"����H��!����r����=�K��*j�!bA7r{܃�V��a�L�/�X��0S`�ת1���~ٜ%7�V���*��q
e6d�j���,���qa��v�����|�(6�h(��>+�b�}����Z�?��	��B%+F���NH*G����(�7aڤ҉�g���l@��%d+%Н}<Q��q�j�h'9�R�w�<���(wW�9�E,DVf-�ľ���hfX���x%��#�?�I�>3�f!q�z-��>���[�&6`���Ϊ2V�0����OSaW�#�(e��;��g�B-] d�ve!X��:m���o`(L��@nѽ9��I2QT2�
�_��RdHᲯ�D���>�~
9ْ� _0�''�Y�o�� 'w��V�K��4|��h��f��Dw�3O�3ڳ�gSvsؙ?qsJ�뀰1��!��
��h�$�l���Y�"�/���k8͢���AQ�q�&�Q�QO�ICty��b4�w<D���&WY�јFҜ+Cm��	xş��l7=�.Z(����J�,	���UN~	�.��i�b����HS����LB�ޢ��z,�q�P^��Q�C����e��7�Gkƒ�6��d����I�Zj1���7R�}i���#�4��Ү?�J=8]�a���_T7�ɵD�p%<"�h=*Vc����˯��������h2Q�x����O���Ԕ?&��"��!��Kٵd#}�T ^t��ɕ'ul r!�VV��i�8�-�+}b���w{�E�#�k�Qj
��K�CA� �dh���D�r�e6����0o]���
̃�2A�6:K�`bQhW7 ��S��jHtlqƋ�t�X'F�ݰ���.ޥ&iN�#[�h�hg�Qӹ���e	�4�xP��LE2����q��B0������G�]�IgS������T���������4��?��5b���؜HB�R�!gf��r����z�Z�ZT#S���
�"=z��Y%^"	�QR9F�}EВċ;�ހ}�nn��u�r���T圣���&]_?����G\R.a�<�d�L�
k��bM�a����l�N��r|BOJ��S�ٺz�ϩТ�UY+�J۱�b99�z��+������|D�ޜ�T�_9�6��/�c~¬����EvO��ۼ�'$r�X�<��p룼@F�v,A��Ʋ-���9���U~�)~�u�@�]���%%H�X	�wy3`�Z؇����^m#��ǡG�ɀr�R�C{����T��3L�v������-���n�8��q?�QB#��!SNZc�?i�� ���q�qn��ϥ���\�]��3��1\��n0?�s�!QLy;g��{e��%L�9�TT����\��n�>-.���Y`�_�u/I)O�J�M�Z�c)a�4~|�ȭ;d ���=1y�㉻Ƴx����l�k|�����g�,W(��s��82M�]^�?�*E�p��[r�Q��:ת�o��R>������w�ce;�v��V`L�{yjd�xѕ�5��y��(L���w��ԝq�(�V�hZ=�{�R�\q#@��#)	�Qy�J�H���s���6o���
�C����(J�33�ݯ���.it��v5�S��2|]��I�}E���.M�9,{�����>�N�+�Yw��f��1�"aK:�|���}i�4�����K{m�-��J�ئW����I�����D�PA�XY�ϱ�U�^�]~�t��D�\̾��AJ������'�]Hي~h'SG�֗����9CG=,�2��D�Gn��x��n�kSP���"�Vә��>��6�y�U�!�n�"��D�g Pp��:�ʿ��r�A��*99ç��_0�����$�?�v;�`z� ~#x��W�DE7D`'�ϯ���C.�a��e�_K�	>O�z��-6%���X��� ζ�C
^�������* ڜ+�-��ӻDҰ��w�@����2+d���{��?i��$@r����)gܿ���T���n�}O4='�Y3�qׯ��SYN���5�����������cu�n�1�[��2u�sx���%Ft�O�0M�5[�(����6_G���Y�j���yg�jr�&Ir���f!������V�,C�����%`��]��&���y/�>�`C��DA0�+�7ǈs���TGy2�]G��1�� �Kst0v$�?��[V�.l	H��84���=���I�k[���(�P�����܋�딲Q���j�;�I(�{7a+0Tlz�nN��f"�DU_�~�nE��]��0�#��ղ\�H@��G8�O��`>�&^�7h�k�[�x�r��w���!����T��c�u:�
�Y"�$��a�gd��c:��J^���s�ԡ����缾�۵�O.rH�*���\��r�.�?:��T�+��+�x�����2�
��*��(	'R���S�[�#9�{1w�3��ɠ�*@����c�e�� 1�M|�Ѩ���G��Z2��x�B�6j�g�=�
������/�$E+����ϼ�1Z�a,��〃	g���f�.�5�'U�*i�7v����5�M�:��P���MJ���fq�[��.,��.|��6�B�[%X�E+����ծ����
��B������)a��ݞ1::��ɘ���\��H����W�P����>��xH�ծ:� ��zJ��ε�Q��-�:T�kT���2T?��[I�6�ad�R�?Pe?��ߢ3�0w��~��:ЧE1&+���t,��V0�c�H����#�}�f�@7f��9�wlSg��1�¼=� ���zV�6�A��Í�/�*A��?�X�6mu"Y�6tH������Q�Z?A�q���r�?XKY��5�@���b.�Cxg)�.
�Bv)��*�6xK�D�K���_�9�*��
 5��XI��x$���@�(�L,�A����ޣX����
����6���ô��/�̃Hr���X;pr�0z�Ƃ�N�]�Z�K*E43����Yct>/��v.}���)�+~Ҹ�%�c�s����H�
����( +��م���8>��{i�/�d��z;����=��K�Y�{��^�d�
����L���AU}�4���-'P`">P}xR�e�����ۃ�Mc#�f�ۖ)���g<�~)��M�љ9f �Dx�p���1]�7X�ё\k+�J�M`�%+ʘ�=�F�����,�2PA�Z�tJpl^�ڸ�8�-�e�d�e��}`m�h�!H
Ż/����5d�������`1W�&����3�( X���LB=�EK|\P�{��R�w�V��륦�c7j��:��lt�L&giݦ̓e~�i&��lJ���mxv� 4m��z�t����_0�����J���̨"��fawg�֏�x�$3Q�Gs�5��Eo=\�Z��������|	p;઀7�iP��t�x6�'�d��hS��Q��É�-�������	Ю=z�6_M����h �X�:b��"�Y��n�(2��RX���:?�ۻ3��.��<�p�C�a#$�v�=�2a��"�b��� 3�*���Ի�%��TW���Ъ�V�9E�Cs�}l�����6��8叴��M_�cP��{�<n�h$(���j�)iJ����QZ�ܫ�dKD
�1n�[Q���Tk,0\m�t��#�NJ{(d�d�Sz�S���*�=�p6!�]�|N�H�U�]1���%u���ᥓ`�9]�E?���wLRYۭ���2�'���
�'�e��3��m���-��u�'S�e��Z��IG|քU��`zi�.م'�����C�M�c5lx!�'p_���՝#'����ȫC2�Χ ������n�f{��6�Fl@5l�Iyl�����L�>yC�[td\4��ԛ��BnQ�F�c� }�.;}&?*_"��<�$AQ�݁jz��$��a�?-�?C|]�D~�&HV�F-�������K���¢�	h˩ �����~�����!
M�PV";����s�@i\܂��؁�sD=@�T� ���hMJ�o�M�ko�uA�
+�t��0R��"����K�s)��c�s��	�)�Y�"�R,�oO��R�����oq�b����L��a�����[X�, ~�	p�J"|�� ��L�Z�S�}Ӹ}-)A��W3�N��;M'��
b�٨����.��IW�e-��G�ځ���j��ܫk{c
�����S��@�����/�yJW�<�z�	e�4o��0@e�au�52���ͥ����.f�<��:}�L�����>FL����k�L8�\
��l���R��nV��u�0�M�刼�Q���.��D��H)al٢��-<W.������	B��㾽ą����-ʥU�j�<k��}/�������3*w#DY/�-�AX�D��Of��&C��-=����|�� ȝ"�/S�֘�FlyӐJ��n�@tH��#FCf-��r���s	���\�آ��N@9���-R�Y�w��'���x7��ڡ����A3T�8Tz�E׃���~L���ϿZ�4x�I\#��\g�.HnLN���hn�G�f�3-�x�q{+04h����?��s�QSQ�M�_�Z'=�鄑D�UVB��>��N#U�@����G�T�N_1	C�����En��;�]�-�XS�_yy_%�EJz'�
���$hV�����J�)�֭���vi�U`ok�"�+h�W˾���&����~��)���������d�:k�Q�������&n/��jɝN"_��Fgϓ8��aܳ��������F&��̠5��Iix��S�áQ݊��P���?�ޠg`e��;4x>9Wx��N>Ķ%y�M�kB�W��O�p}aA�C��Xk�0zr�c��[}���쫸V�Zv� ^��9)x��wV���ŵ:,a�ɮA���5@�~L��ŧ�U&�$�D(*��v(`��g��p'�!/�
&�k�bl�i�+ro���E^�
6Q��к_׹蝮!��i̋����n�ك*L��3�凟�\[*5m.���o��N��N�S#$!n��>�c~�?�<[:� ���=[�7i�nbAfd#U��k�v_�M���E/N1��� �*喋������j�ԭo������Vj?���\�>��y�C�J��Y�	��oA�w�d�k6K <x4f�V>�(��J�{��<��ܤ���YBȁr1"����`� �/�3�Liކ�H�P<���BX3+c"�Gd
�j����y��$7�ܧ�k메/��{}$�3�;�/;^~"�NL�R:�:�h��,�3d�x	��>'Y�07���v\�Ȳ�l�v, N���0F��M��O�p�f]���3��E�������>_v�D�
߿�էr���н����g5�`�o��C)]t ��=�K�?� (A�&��-�͸<�2�ͨE��>��X�m�z"���K��}�^���_WNx�����m��j�m�_�]���V]e0���z�O*	@��q1>#)���-�7���5��dG�ʝ��Ϊ[D�#S�ԥ�\[j��g�Ȣ���e�r�OFz�����L���WOJǼD-?���V�uD�!��ir��&ϑ�y���sY�Z�^��&���⟇lr�`c�1c��|۶�Q��C���/����܏�O}�F�}���Ͼx�ξ�=�/��ШWIn�B�f��܉Q�k��]�Ţ���SP��i�$�?QJ��Ю��h=�ϭ��P ���F��2�~���ô����C�<�ٽ�l� �!nԌ3���$��%su��v<�����K#r1�H�B`2�6�\�.l��Ch���B��{�Ep�l�BZ^�*߾Ё���>$k�)��ڜKp�@�l��]�%���K�V�X����]kZ7-4��O��|Ħ	D28ײ�v��h���#��S��κ]O쁪H�ǿڽx��}�{9����úD�N$�r�ZB�|s��8��yz�`��"���\�'H�/��-*�l�tY�iȼ���^�Ɲ e�Z.N����ԓ&ǋ�]
����r{��ЍG���~�n�&�J1U��@�*�m��I����X�~<l.��*%����|���Ii8�������jJ��Q6fuh�ܕ$������{L�3K���iQ`Jo�cQ#��f�*��;�q��5\�_r۱2���i��Ӷ�rr|�m��N:D�/C�x�%�R3��=Qr1�mE����kɢ/�X#��Q+�&�0s��?�tIˢ�􇞉p�*�+�_D�I��so�8{�J��̑+)��FJ3�~A�`��<��d���ծxV&�?��X&�L�,�D4i��X��i怉�"�)�Pk�1��8����}��L�b�1�6z��6$�d�`|)��lq��c�����=��u,������=.cRjO��w��I�5�W��pp��r��/יxv�����g�Mέ�e�J�݉j�2t����%�����?D�'���t+���kg��)g����G������l��M�QT-4�����X��3Ȅ�ٓyاB	gy'N���-ٔ?�;71��SRU,����'���5Y��i�����f4 gm���:�̗�����=��j<�d���[�p2?a�H-�b.1Vb��n�fB�K�o�?|X�:��.W���Y Nc��5��"�G�p@52mQE]�]|�
�}r�N��v��dm��9�5�M�U�'�F��y���@ag��E Q��r;γP
@i�.b.�]���Y���F�2�|��j����������v���i�Ki�U!�n�W�zQ��n���M�:9Ѳ��m@��'��f���`6|h|��B?�0ܻ�X6��	��(��e_�����4��x�d��3�J�/N��{�n]���gn��5Wղ�����W�8���]�Rdp��m����ǵy@��k:��54���B��ӿVݷ���#�Lm�y� �ّ.m�%�;�[u�Jb)��/Y@L<(z>��A�{�hȋ�[��`��{$ �!��Ǡtsqn�z���l�ļSf���=pxJGf��R���0��֞�x��3��Cȱ���� �J)��¢)ɇ7�7#B4CA����L�X'E=k=���Jf��f>F�g����4�8�9��aId8�2����Ď*�G-ًt��trʰ
qHI���F��k�'tv���s�9�)2f���D濢�5����\VuE	���vF�c��{b��$��3�IF��;� D�f�Ui���.(*X�+�-GP�8�}��.&U���Y�L�A��r��x�<�ɸY���iARSXR� �8�0U���6���'<q>9��a6��%K����:��ҟcM������q��s1!��,,��.�e�r����6G*��Y���p ����U(zjx�E�vDe��l�,:uػ�c���@�@,d��@���� �O�Jl�\���E��%"&���tX�^��ڬPLf
�s'�� ևR�W�)!jCP@����gdI�7cV�c���}'u&��>#���󰶍{f�gS��I�=�KFFLik��J� �Un�2��u�V�M���	�?�\�jE��z2m����6�q����>R&�����R6��O�L��^ �W��u,h�؅�O�����5�Ke�Lzl\���p1�����O���*y�X�ӏ-h.� 5�*^��D'�4��h���o�N����R����	������1(:#O��uĸ����r-n�m�ڠ��ƍ�hy�URGpQК���#�32�w��@b�V�!�����ޗ�����h�͍9,�T�6D�q8F�s�fN�e���($F1���:^�.���tԚ�e��+����WFW�iW���8�V%��48u���W��R����y���}J<p͹��2���2��Wg�v3-��`H��,�2�0��<#�bk�G�"e�{�Nw���W6.�h8i8�-���ZH�/L-*C��3�V/��1��}���Or���ӧN���n2t���7-5�G�c�1/�4_E�������U��$�ܟ����4��:4�0d_��GaןZ���yc��:��|��Z��Iǐ�O䬸��D������,L��C`��x�ē�6L%�x ��j��T '���C��i�^�`�)���ҩ_`i3N�d�,��;V�"k��r��Xt�S�/E�i��e�Ƒ���;\��ZA��佱��ꢙ-6��A��E@8B��k�/t���ӤG�JS�_�A*�����Y;T2U��Դ�y�=9�O�n}\onG��.��٫r�_%G�U�K�9 pbn���R��)�1,17�z�'s,#�(��=-��f5GK�|�H��n㊔�Ι�*�R�O���ҫz����J@ cu�~�;|r�R���~�S�Ber�7 H��1�ޡ"��@P�L>���5���5�����|q?��v��fǪp7�~3A�%�\��n�S�n%���e[�>Ɖ��4�2�E��ug�x$0�jP��R�{��#�b�N%����6�� >�ھ��'����VF��P������I(�������(4�ee�źǕ/����peǭ㗲UjـrA���W�}(��lM�C�"X���D/M��=�r� �hM�	��,
�[��P3aa���^��� ��5ҋ�I��-�ֹR�	};x(a>cI���S��|d�O��jU$�a��|'T>m���QFJ:��0�a	�?&ĒAu��01��K�J�_�\��%t�A��3��&,����f�$���#�<���Z7�p�le�keM��AČcLk�*�Q�hf�y���Yڤ6	v���*�~H�N��s�8G�]v�[ gG��P�(��1k��J���8к��DJ�q� �շ�qC6��M�hx/����2���r2�X2ex�J���h�]��z7�Y��f&�(��(�#�j|�ݣ��&͂���Ȣ�bDDl��H�*A̍ʙ�/F�\C���%��D7ۦ�R��+�UJo;ݖ %��F�������R����V�]�PY��S}�(�|SJ*�] ��-��Y��݀m�s���(8�����V�d�k��b#Ri��wS6\ov�K��q88᧒:�\���6Dݘ�5��W�;y�Q/c],���\5���|�f�����i�{]�&�Q�9�C/ǦR����~�3���Ц��w�˽�D,�r%qiS����R��:�uyM�m�9�a��P��T��'����󨈒���#_�6n��6��8�����˴���$���D<�� )�����(��>��p�A|2�k�k�@\T���:V�7�#�zOG��4��,�c���s�1g�,%�N�E�Nt�����Y�0�՚���b���ns�P�B���"��R߈�6��޽pj9w��t��wT$��f}g��k�[��^�ؓT��4mM��Hղ�SrN��M�R6D盡���M�* ńo�Qm�Ałj�	��O��g��v���J���r��y@�{��zk�l�B%�Fgn.�Pj�Ur�,s����]XBU)Q��}B/Q��NM��/����k-ӱ� �$��.�Ԗ�:�^Է��E���p$t]�ص|���<:ֵ<[	�`U�<k(}��du��%��`�j�Yc�Q�*�ރr������\g��i�Vfg����-��i�f�qY��@$�[~����ׂ"�C��u��C0�5ݚp/�ƈ�f��6��jZ �	v�a7����TWZ�$�ؐ��aQk����+�-�L	�d��*��v�p �	E�Sg���R�bN�5��[�*3����V	a�/k��l8R�lUM�~Z�MGK��<�0���}5e5�R�o���9@�/���:B�L���:�$�K ʱ b� g�RU!��%���V�Ӵ��k�@�)�OT�96�1��m|�픔�GҒ�^����?�gĀչG���,�ƈu�XH����ՠ�s�X%��kP���B<�Hl�g�Jx��X�[�����;ڜ)4��q�^`l�^vʽ��	�;��P�k�Ί��7rY�\�`9n+�����e@��tO�Ԍ0�r�yg>��4~�2И]'����cJC�:"��W�����N�rȋN����-/��b��������p�z�&�[���] Q�)�5�V�Q��QF�F���a��tw��$0�]E�W�de*>�0���r�1��5�f�M�ꮄ^�]�@�e����>BjB5)�Qm�$`I<HW��u�F;�;���"��*�|���k#)ʐ�2<t��F!� 0T�ul��v��7�D��}�)�ǖ���ۭߖ�6�{չt_��vl���	���s���:V1��Ph�~���h'����#����ΫvKp���F��:ȄHL:��4ov���'��/A�����&��E����1e���(gm��@9����_��Eb$�}7ؒFWbfo��n��P�햬˴�j9�Gy=m8�=|�^��f��7s.��F�ACP��.ec���u8�R��*���ȸ��	�{�K �-�A�s��)�F����U8F�x�#.�W��;���T%N��:(+}ۏ��cӈ/Я�'4������eE�M�q?�5�	H&��Z�UT�1�4�rÙ^��;�2a3adϵ�z��(��zS�Eq�WH��O�1aAͮc9M�i"�K�7>].Q+?]nŞU�6=�L���sJw�!l4��`e�����Vp�! ��bd��5T�(��[x	���A�C����GIT�B�O��,T'K׭�}��R5)�;���}к�.f��C�#���Va��8��@)w������%��҉UH͟_�u�3X��Kh�A���azsGs���p���^���������#��3�r{�~�\1k,�W�&J5Т�|,3gҵq[u����
��j�����?�+�:��w󁑿Z:>{3���r(q����)��A=+�k)����.�!+(���7A3�i�!����Z���������;X��������I���}��V�(W4i�o�h="�Zo�@m��(2~H�v��kK �rՠ����%�a�Ps�dǀ��RjU�T�q�^��\���Ʉf������F�T�v()�\u@LK��fo��6���K���z��p��S����$����hEsgV� xve0�\�3�RZ��g�u�B+yc��U�l��ڱ0��:���n���q�9����Wʽq����p���1�Wnt�FF%p3��K��ڶ�p8�0@PV:!�h��|)e�m��UTr2�[X6Z��N��zb]�x�tw���$����B3��;z�U���ʡ�FY"�L�{�홄���j�b���4%�]���D�	MU"���.1�\���)�����x������Rp"-��0��de�ѣRA��ޕ~o `�7k�(e�Ӥ�,�=�^�M�w]CM�w���w����3�c�q���O��-b����B���8M^�k�����?��~�ڋw��~�@
e�iPI7G:��w̠!� �e$|ۣ���%gG,�����dm*+�V5�D5cI�%�.��4�]?�LY4��ump�����/
ˤ��+�at��!�Ŧ�J����BV��5(�G�O���W�z<zr`+:�Q�Q�ࡧ�-��
���<>=<j�\'k�w�r��$��z����;��o��u�|�/��G��ߠ�OD<]��~�r���	�{�"i��4��L�6�E�b'��I>lکD�뎇�7@&���l�-ka��f3��¸('��u�� ����{�� ��Yvy��N�?.�o�gr��%OǑ}�2'��$�W���R8�;�9�z��ƻ�i��%/0�PB?�d�,}\�(��qB6+�g	���H���z�'�S���#�ߥ��o���r��ʲU�})i�H��0���Gc¯j��"�IR�����f�j�����HАv}�4��c�-���ޓ����� H��*E�=*
�+',�������ARK%ψ��Gv���L�>���ǣE���u5-dr��b��	�Tlnc��q�J|k~f�sӎ1��\U��O�c��3�iG�q�1+�~�\�4�oVtC�A:D%�7��D��g��l��1��C��j�ȝ��`���@�-��H��G�1�Y���뜦�u}P5W��R<�;S�N?>d"�qW�Я6JV<wR��L �$���	c�-67pu���� ��Y�Fz�*0]	]��no%N"�.~���Ll�l��Ĥ��Z��<<��l�V��fcU޿��s�9����q�"<�g4c�b�"�U^��5�g�՝ٺ�S�H٣>�k�g¢�;P-Ҩ�c��4O�&JP����"z��{F����Ջ����B����u�mX�%H3}s?94Q�ꎦ�8����;Hj�B�p��S���1�"���'C|�YB�������YޛD�$���;�k��b�%�YN�W��X��y ��`:���>e������tg��b��b��k ���#0[�����x�	�[C�b/�p���׼���s��c���3�5���mp'݈)�X΍�X�����P('��9]�{�q��yu�J0^�L#�0a�k�v��3T����x}��(`mqx��Er�*\RQ�h|N��F����Ύ��4_�wb���~4�"?f5h,����,௑� B���2�#���B����ѓ�13a�:�Fj���u��<fEfY�����&����c,MK7-x�r�rvQg�6���dV���·��,��M����_A����N��2���m��B�3���U��ܻ�;���ri�cM��Je���s��ד�U����m�&��G6*OEwE����A(��E����L6�� %�8��	���x(���Е��l:��U���S���|��8<jJ˭�R;�����wqh�0��1S�p�0~���B�LI0�>O	&wib��"�����t	�H�Dw�9��N]���F����3ڰ�i��،�T�2�b��4L���E���"[�e��l���9ɟ]�����n����[��;� 0�s�EE��-l�Ƞa��I�}u͒j/��w�X3S�4Jb �ӭ���Ho99B�;�,�08�Ⱥ^!��O�_�aC)YF����lF�	@<�j�Ew?z��f�r�|��ͤ_�P�/IKًX
��L�xN�LT��bWe5A)1��u=}�}�jK����i����x�#W����	�����_2Q�1�	-�I���`t�`vT��~��r�}L���5��c��Ph!�?cM{G�,!$���s�T����*#"ϟV�X8�.��SI
��HP�� �C��c+���OA\��V�ߞ��%�)��\5I5ͻH��l�+�eu��-�JTY�Nm����]�Z��fX��;�����kn/���zk�N�yNsֹ2{��E.�Yʼ��>y>���g�>9ĕ���*��ڞ�s�M����Ć՝��?�߂��~�oL%0O��w[�]�j�Ǭ��賡�f���`�%!��zg�2��@�Q+��/3��T>d��O��K~�y�R1��f�0B��?;���������m�?p�#�K|�T�hb:9! ��J��ֳР�\����Z��6x��m�na��7|#���<0�N�Z;Uh�n��X�1���'ރ	q��:�"Uz��������z�<�6�#�u2�t��m�¹�I�Jj�OT[.dq�e��b��HU�30��f�[��nV�j�ڷ��H�@��	��{f�"�HM����Lw�Lc_���+_�8HBK�3��[�K���5�$w;�2�rnԇ=J��?D��I�,x�����$x1@��;�-������(�疩��a������)Q�z�+��K$�$��� �Ӓ�jY��}p^w��Vt�����$*�q?@��,�p"X����{�O�޺	��w�،�G����C�e�u#|q�\8w�����Pʩ��U�]�[��;�ͪ4/���"�c�������\	]�=C�Q��L���ׅ.4#���-����iq�13%��d�$�ϵ��*�!���Ҍ|����柹X��Y�_� JʘQ���ү���=2�K
�1T�_�dP��,ս
��Cd�r�z��J����m/�P��Jvq6w�0H!���
%l*�}Я��%��L�f]�A
�ĢY��,2+,,�tjF2�{�[�!{�w\��Y��թ��X�A�*��؀j�E�`K�~�Gl o�*�B�"���~^��";#���<l�e�@F(���Pu��1�y9��8U�E�͚���1��|	���Uj����6�Y�#Wb2V.�6�<zF&۔.��T���O�^�
�w鸧b!T<�XԴ���ҁY�zCr���O���\EB�F��<�����"�ʔ�[?��i�Q?D�Y��ux�ϝ!zG	�D.Lw@��4#�t$X�p�?���5�/+<^�E�B�1l��M��j�ˁ��~\�;�xJ���M�)�;�Z5H���Q��}?�wS�9�_O4�.��IOkblj}rjy�=�����q$�U�Z>͚)���Íe�����2�2���\��[_ ��~Rg����_�����yB��t�3�����k�3��:.i�<]��f`�i���/�JM�����-ff3��+	<�2~��v=?���em�����m�&�q��fE�q�]_x$�A���2���իV|[��]B:ۊ�.d�"̹!C%HzːM@vf
�[���NKx�g�M���K��w4Hbb�d�em����#ݹ>�!چ��<�$8�{�¤�(�����_K�pn4�74q	(��=J�%-j.K�k��{��z��[��(��9Ƞ�1Y�=ۜ�	����XU1�����&)�ՑS��o������=9�Q<T��(���>���|�8E�p�#���#��h�$!��R����_OA�r��ǒ�; �6@�X�Q���咛B[߁R�#F�hhQ� ؏�fz����`�a�֨9�i�z��Z�w}��c{b;|�c4'4���}����Kq�!G�I��p0+S�c��7�,+�O(��r�ڂ�@5��P�V�o���C�fF#�Ǉ��Nv�r��C��q��p�|�A����� �#o�R_���:G���;?m�D&�Fn2�I@1���O����kc�O���S�*�<��z��MnWK�k_�5���u@.���%D�5&7��9W���� ~>p:S�M��tj��������{p/�1	1��yL5�TϷ]~�X�S�P;xdH�P{C���&���]�����CCP*��r�7Jb�^��	?�����0�b=���D;Q^�C�0�����PEi �ᅹo�4��-C��N�����&����[��S�8��kœ�Z�Y[m���gηC��d��(?�X�<H̾�������1�}���o;���֢���� �Μ$:�_b��E8�X�����9���M��B��O
��81mF�puZ�V8~��M�=
@��K~�Ύ(�_"��3K����3)-��V�n�,T�HNe	5������o��(A����k�L�,��1$=�
�$1���n��-G�niu��/(n��J��y�A	��m����=��M鵿F3sZ�U�{�٢��翭��ʗ��-���'-�1r��=��~�vE剦���y*��(�X�k�xf{�Vu������ƅ�.�3B�9��Qj�?)��>�xss봠'�_�4�Bld��W-�Qt�ț��xO�G���ݰ��xi-_���f�cz��T(����/_�c&ّ!��"�S�6u��Cd^@�P�uK�1���Q�	�yl�mKx��;(��,�JÒ�>����7Iu���m/� )�Z�����*2X��$��ung^�;:����b7���!*����ՠ�����ܳ�_[�0iia`A����KID6�H3�zyͬ�tMS���q$1@�Qm��p{/���0jI�-������&�����<6��� ��"��Ϡg�|H�� p����[�Wh��L�ƂEv��� �}�+�wt�1-���n"��a��4��;�Na�8�R��`�����P��y18�X��5�	}��͘8w :�� ���fN�G@}e������+� �2��.?��������
#uIK���B��A~u��f4�U�$0��Ԯ�D�n��s% �󷣷7�4Z�q�J�̤	�%P���:���)���P���4�z�~�wX!!b�!����@�CP��W�@�8��WR���[�e&�	��,�۬wSf��o�@���e�e~��r#=���A�uXFA��{m�l��	��q��6\=���A�I=zυWAఞw�Z_N�k8A)��
��7E�o�sE�^����vD5w��zX^ ��$n�
/SӒUX��� ��#�z�8 ���̠ei�Xz��i��O�-Z,$G sJѽ��9�k{��#�_��a��l8�v��]�4�n�U��r��"8�4` "�%�� ��\���ℚ@"�_\e�%=^d��z�%U����@�B�[T��gAD=1��W�B�;閙)p�~��e��(�e����P��g�v=�N �Q�h�m�:is�V���</�Hs�,��멻_�d{�$�1�3�@�]����X��G�l��x����(�4��Bnmĺj�M�\�L���� �R�����U(�V'UՁaT��Ոl�q��[UM*x�fF%���'++��T���_~��H7�{��i�{H���}_�V���\��1�}�]���g����.�j�Qmm�WL��
x�8���J����|�OoeR��_���+�*�[U΃T8�;�A4�2Ra�]��m�W�罼<5�'�\�\������K�a4��!~�Ȍ�$j׽g�1@0�	�z�/l�����'Xګ�1��h������,8����r(₡�Ue��HL��r����7��b���9��V[�$5�OӔ��E�;n��7#1G0� ��a����DW|�bk2�`�N��[�}�(����R�W9r��/#7Z�g9�y�5��!�"��,M���fɁJ�+2��˟T&��).s�=�۰+]zY�_����Q����4漐o�i*�Ы�ʵ|���0 #6��.94$�
]�����4\�����x5���s��RfV�]��ؿ[��=7}Z��q��9���9��o�Ȳ�ϐ������$�$xV��b'�1�9�Y�u9┞F<�����@v�T\y0�Rvx�wPq�vA��pI��"}B�6x��.��b����b M����J�,ӯ?����NMd�����O� `G��L�JM^b��R�-��,w��4q�ژ=��� N)��z{Z��F�x�I��Z��"uk��2�o(�ȱ}�8k!����
�$@eV�ȁ ���>R�+T�`�)��m�g���j#��]���7�y�3f�q�#������0�m�Myu�a��)��e~�Y�eH�L����!�p����ݾ����N{䍅�he)(��i�՜G��?�4������4n���p��C���� ���	0��D�<n��C�ĕ)�:���2����RM��A6��+s^��m�z[j���?�S��EfUr��2��-�
�d� �j�G}�`�NuZ�
���&m��l���Y�x�F¼ST<���7���Z�ߛ��!`�ǭ+�8Ol+H����������/��[IK�4��(�9.�3���)(�e3�S�!F���|�g'-Uo]*8��"��qu�-E[�v,м,L2�H���8� �=G�|3���>�yd�
Ȧ{�J�ӽ���W���ꨣd�P�l�ӏ�w�~I���!�&�}�z$/mI�	��Xr6	;7@࿨���9 �����
ms,�pxy91�r']�����
�Ő��E=�i� �k}=}��;T[���Jo�����.�d�$E�4?-�4����N��4�Ro���{"�Ŀ΂1SX,�-�\����3��16�"�-iْ��w��N(�{@��Fdܮ8��ȳ���e|=Lȁ#+�/�%sі��u(���?6�8'[5�=+Awj'C0b��D�hP՝�nx(rv���6��>[،�ܬ��w ,��=(">:��ڿsXdt��{D0у\�T<�Lŋ���Hc%�_pLDq���/��]S��*��h�����0����6 �e1�AU`Q̈́uk:'p���!k*1ӧ���h�M�!���u��@���=�F\�D�+rt�!;�m�&#�<=���CwdȎ�\Yo��[5���!|,���߬鳱�����ŧ&�A$T�u2]GJ���� �8}̉!h�B�2�S�j%_o���݆�����y�1â�BM��ú������.C������@Ӫ!�����t��P��0I����en��]��}]@	L�W��7i�<�Ul�`l#���˹j��/+��-G����a&��گx�%͓�n�`N�_�x��t��.�T��&Wh�.?|<v%��18�4�9b�zZ�qQs��:�Ċ�HȀQ�B���Qڹ�U���,�+�[��,^�#Mx�I��o�&�đ�5�K�� %cT*�>����������~Ѳ�/7*]���|�Lbmwv�^4k�3Y-bzW��t]�b�ުh��tF��$�5.lWU�9>�6B����V*s���5��������b?b/�s�뜦������]Jy������K�"����`�����b�`�wP� K�$��5�
Bas��t;��K5���
���g��?.����g�pʗ�!�_����o���v��D��
s���?
_\�a��R����40��q��ϧ"���b��β]xL��ԭ�*��+#=]-d��)reڝ}ڙ$M��P����n@p����#���W|s���t��do�gF&�8�>B�E�
0���,@{G���$�e� y9M�(�7�q
���H�̩�.^�ā��<�\�RH��H��B�VU�D���5qjr��WG$����K���u�T%�R�p��үA�.Ⱦ�!��8�qA�kN֏"
Q�>�����-��(\�08I^R���9�fͳ�5��L�̴���i�P����0�!�����3	�!"� @d�!�sBt놁�a��)��YP��H�9:?s���<-�d7�2wR��j�hD�C6��r�7�u�N�L��@τ��'�m�Q^��Y����⭹q�P� � k_C|{ԷOv8x�*�|)��`��4�`�8ƒ���-�@�W,�o�9���K�ϫ#�g�s��r�� 1'@A!·j�k^Yn�����a|'�FH|��ɔ
p�|���h���0�[יMr�! �~�P�_錪���+�C�Vֻ6L-.P��{ZO
�aTt�$a�k2���̜=�����B\��,�$�CJ�Q��	m�}������ay����4x Ih��%G�Qp�VK�����g5��X'֤���7��sڄ.f�x-��H�]7�L�����A��A6��H
�dsI��P[yՇoȪ,�����ll�	��`�UD��O����Ž�iw���)jJ;�u\x��4V��}G}<ݲu�en#����-IC!5�9�d~�ZBu��6����u2+Uyv9�s����?B����G#V�<��z5��wxd3��1V��g��JN�ñ�ɖY`������3 ��\�F Q��ڹ���c*�J�SDU��k�C��+D���5��o��h����Ziy�-G-!���������q�kY���{�O�$�����u��j�W� �ٔ��	nAsES�����/Ǧ�e#�!�EA�=��	j/�-�����ƅ$�+S�4����EĶg��t�g��~�:ai����S�#���L,y�ȲN�4����	c�I�c�v݁�}&�]��A�i���h��	��
��� q���4a�c�H3�3x�b�X\Y1ɛ�	���a����HX�	�"�c���u�k� ��p�u�=Nc�p}��y���<�����{���m%����mz�(B$��t����X�	.���ra�w�ַ�t����������H��B�d�"l�~�mb}!��;(�������i�s�����H	��G]v�����P]vK�E�N_@��'P�2j�$����_�?�7�<�ܨϜ���� >R��jLO�G�c����0��a�C�.��$5�rc�#Μs�\��F]�Vu�����Z�o�%ErZ�nJ~�~~��>꒙k���@`�xď3��q�fJ�[P��'�`'����	&�����>c�ڻ+�L�ˌ����GM\�!�q�h�_�y0�
W����-���(ۙA���7Q������j4��d���@�F�.z��s)�ݲ�sz�R���w�-�mO��e��^>��o�Q�lCMVz���P�c��7+�ҟ�k��sjT��H��Y�"N(���Լ��O,B6����U~����n��4�i���eC����@��b�y�>����t��t��}J�a@6��2mVsì���P��+O��&�NR��+��=ӱœd�������j��u:87�����a����l��&�\�G�h8���8K
�v�Z����>���4���n��=�-z (Q�vg3H4'\��O�d���Y�=��5�S]��lt;��/y#���x����IOJ�]�~����1�7Rz�V<3��g; `h�iP����n^s��v�����_1HC�bp��S��e�ۼL��*�_�q��|��v�>�È��oU��`�f�¼��F�[y�	��=j�52��	�
�jQߌ��B��m\�ur���RC�����zm/ϰ�j���r�7�_P������ް��.��w��e��o}����j��=�K�NJ��'Sm�ܫ��r=�������NM�c��cRq%,7fi��Da���j�O��B��Բt����w������6�-�m�?����'�~��R<�y�����8]:7��F��۶��(mP�9�2��D�Xab�ۛ�Ŀ���iH����#�,�ıJ�5֙�G��p��$�/ڸ*�Υ��h�k�����hCXs������ c�� �e�Y`�e{�#3��o�����E,f���_����4[JU
4DJ8�ފ���Q y�l�@<�]����5��z.>��C����9�`ct�e|��Da糿QM㧮�îό�=R��q�N��� a4��ʯ3 ұ�[9Cn&G~_��bo$��bi��.��������1*Ξ$�C��%1�R�@�ӧ+�G���g�@g��o�gmѭ2��*z3	�CIsN�C�W:12& ��ߦJ��!:�3a8]l��\+X��ȵjsӬ��X��`������:��4�w�>��=L:W�·&Eajsѓ��d�@���9�^*�ia]%����j'�ys��.벤��� �����7��f*jE;C�/������_��t�ɜu�L:���& 	�q���ZO���eF�.���9.��k�JǔЬ��Qs^��P�X�Z'
RL�M�hб�=5A�hf/�ڤ��(�<k�����+Q��;n�m�zF��/��À�8I�ъT����A�H��D6l��o�9�X�3�w��~�_q��v����;@�;�vu��
���ȏ��Cធ��M厫�M����)�ֺ,�u�Pւ����fi~�[R_�F����;Y
��Bc?�oI�)a�w��	��oG`&c�zij��dv�z����8x����d���Z�\{�{�X9SLQn�_&���Q]j��/O[N��TlV��
���I�QJk����(�^�>J4�����EFoj�ϕ��.�����᝾�P��Z�}���maL&ڕ�̛F%�60��(�P%���'���o^*.m�pIQ���^%��p�NR&ϩ5���x��ƴ�n�:LQ��XX�drk���z�vy{���%�``W3k�>����ە�9b_�O����^v�n��7;�D�.���,���	��K,�0��sU-�A�V�'��W
3��&�7Nؕ�h�
��إݤ`�4����e�/�:��T���v���3���$q��� {˘�`r#��q2��N"��,�P:�x��)K��'����Z�q�+�J�"����;�H��rf�f�n�{�G�O����p@W�C������~�y˕+�h��V�9Y�}��f�}�g���͙4h�e��p�1^A�]fP�� W`*#m�*h��H�,��N�]�
�-� ���Cҵ2�{����-8�7��p��(��)�P��U�[��oxuYy8է� R�n�`\�|L�*}���l��m#�l[��)���i��5�(Tgz�Mj��g�4�@H����FQy���'`3��e�|Y�0LatU���亂�~�>oif#&ÄYcԙ�֜���O�O�Er	�H#�.���l�%lW:�S%������DMx6i�~r%�R��skR)��,���y�"��N���*0�(�"A(em����RF��.d�,�̠�M�o�䟚�	�SG�o�m+P��xk7m�ji�Dג�Y"w�^�N�M�}稬��*vk��y>�͸)��.�J�+�I��Z
�*0�ET����OE3]"�3&�y�]�NeQ�3u�upfl6��_eX�,ň{���'�ʦ4�w*��o�u�cEZN�T!���9Z��\̿
hN�[�1G�C~I�ͺ�r�~غ!���:m��a�g �{.�!�E����3��փ�*'�~U�B 8�@O�J�����o~��+�/���;��m=�7�  �˪��R�t�A���}u:�#�Ju���H+��V�}4EVW:e��0�0�~6� rz�d-j�U�� �qf��̚���w.�먇�nie�.n�[�R�xa��UD<�*97�	���$e�����t��������x�Y��θA��q�w��΄x��P���gB���Ⅼ���Q��*g���a�M{���[h^�������� n>p� �B��\y�d�yG�@W����+">-bVJ)U��
�^�Sq��ԫb)4.���E�ޫvz�f�h�yP#�#�ޣ�c�ǰN�Uj���:2���Z:�ӄYY�d?�IG�82�O�ɢ΀�<��Wf١<Zn�QI��:Ռ\~/������w\����}��rM��X�	{P��=*
tz��M�R��eO�g��M�"k��������K`�:X�����P:%��͙���7��@�5�6� ��R��r_�0�sN�������b���E��C�$qد8�y�#`������{GGwt��?��+��?�a/�P�fjڃ�{p���h��yZ��e0X0e^���Ӣ<䥩gSAƁ��xֿɌ榬m���Z�uM}Μ"�)�a
*D�u�;�+�Ԍ�
��w����a�D�0E)�ڲ�H�yɎV,�'�@�?�W�v	�C�j�x��[#Xf$A/��n�
�b�߯�u�����˄��;CF���3�W*�)�d�z�'vB�X'dIûE��߮y�2����3-�w1<��l��{��'K5�y�YV�쐒��v�R�.��{�l��9)��d�$�ܿ0mƩ&��-E�O����ʄx�;����,S6E�̳*T7�|h94��o���P����P�9�Au��2�K}�Q�as���&c�'m_,ɺ:�6a�D��&�(Z�Yx�w�@^��tw���Zo~��R��N�,&����pu�#(q�Ȱ#s��`6�2�Y4e�#�����p���+��t�Ct@�f:ðDLseB�<.���C����.y���rT�BV��DZKx*L����2�Bߪ}��MA�9���;X �I�d��Z�F� �e�0*���=��#�/���o��K����jaа3���*� ���^ת�K�����V`�_M:�j�p2��-�.�7�_�.��n�@�(�b�1� ��TmN�H)�>1�䄇�~���硧� {�E�>m<���:w*��h�� /}��,/V������Yg��4�U����t�(�T^�̅ *w�Ы�Ѫ��d��ԝ; �_�f�}���)^v>��t`g���lZ=�,N�V��z�pf6rm@M����gd	𴙬����� ��Z��F_����t_"��ElR4L���	e��oK�J��i��/�t!��!.�fŃ�<(^��p��0>e�ii�q���8�s����l��=�<�1�g�.=�'��������n�	���i2n�]���c�����&&�@��7'�~���؃,�>oqJ�=�rM�豕��F�^�p��vB�C4���U��N�q6����f7?x[6v������i ���1�7��M<4>��х�#X��3�ڔ�?8�%�����eǅ��v���Y�t};��:��(>�1U��.z����B�A�4�[:Ή�"d{��U���A#'Y5���.�2��Om��%�E�d���*w��x�z���3����~Ѷ�e�>��q�\�<�����-Y��.";�GYXU��*���s'�3�;��_y��9�)s�Ypj�����i�>gi��uE[�:����2~k�ZS�e�Y4Ŋ�K�/��#IΥ+��?	X����N�iXʵ5g��� dȫ�����?٣@��ts��xC�T�)�ݯ')mg��R�8d�'�%��#īAu�I}>�*�m���xKM[�T�"S�q�8����96�xg�7s#T�Kc|��!�d~�;���|>�M��NE�`�v܈Ο����l�7@Zpz��o�.He�w\�Ұv9��M��7�4(��آ���h�_�r�vk�;�n��(U�Y�v%���ǡS<�c)�Nļ�ΰ��/p�����%3#8���O~?wW�'u���0We@�_q�ʆ�K�(���Ff	�H�T�`+t�c���r�426tK)P����r��D��6�=�2��٢� :�,�az�ZFҽ�g=�0��ck&͍��]�M��� ��.�s��G��L�r[1����uc��z�z�חi�+}����'���k����} �����F����7�i#�c6Y�����*�Zh:z���dR<mح�W�%
��E1b�{���W�%����m�;))��UN�{P�|.��9���n��PF�}�N�J�w�U�7ߞ̳	F���gE�}��^0j�ބ��EVy�B����T����w"��U�+8�H�r7���솓����T�K�E�*g��MO&^a,6�b7-R!�2��06���[����x$ �yu�4�ԓ%=�c9���6Ո��p0t�^Ϫ��W߱׀�66:�oeF��?��\�:g(Er�XPE�c?��)^�ީ�Q�t ]�W+�H�\����L:6v@��-ҠSN�L�H,�,�9����3�b����^��9~�������z1ࠔdw�l�G|;55-�d�qG:�"n��1����<K�Vo��i11x/L2���M
gC/�!�:���!�������J'5�:�N�'J}C�-�=���w�@�=LHε�
s�d���Ҫ.�-���R��,���$2�ʤ�EF2fN��dt�T�1����F�a1��Kz���kF1���i�n��,1=�h�o����~ىD��
�8�
"�iha,���Ttwc����f���o�x�:	��÷H3G�[�p3���b�g�H��6un��>�`u���ǖ0���=���E>�- KVe��̇�m;�r_���K!5s�u��7�&�[bE��)����� �?��|�WЁ鞣ˬ.Y�4�[��77�'�p�i�xc��6.�:�i�����>�n3�������˜�
��y����� �����P��kͷP��Z�uTwd����Z����}Sp��\.�~ Ǭ�/��~�V]�]�p�����8�N���Z���u�g�ZN����K�`���e�B��5D�q)�u����MU[��hw�p
��x�lbe���r�j�g��K�|��\V��$LQ����,���������뎇�(��B��G�ELY���ID�����A��NZ�Zӵ �k��y2��*�w��Y�Tέ-K��jp�٪����J[Rݟ�hW:��"x������$��66�W����V�9%���|�&,C��6jI��(C�6��k���ۧ�B	&��U��xYH�exbtY���;iw��x|CO�T�v,�]9�"��A�L��ݾ����h���:�I�8ˋ�r	�+rXx	`0� uj�('m�`���a.'F��n�o.���)q�L+U";�Է2"(��l����m*ꄅ>��s��z)�y� H���9��u3��1��Pn\�����GsM������$#�����]�q_��9]�>!�j6�Cm;ާu #���������2y��c�MgJ���9�ڗ�����N���|��aInkT������f��pk$?�emÞ:�s���4���m ��*d�!n���o��otT�N�f��P_Ň��QD#ʳ�3�����A�: ����R�����`�$�&X�v<x�S��ǃ9w
 �Ｑ��.�[?R"��*���+,��(�o�.�D"�6|�A[m�?���VO��m�<]as���i����^Zd_-{��G����m��VD˟C�6-<�" �CQ@��:9�4��e_�V#8U��
5�k�
ձ"F�J	���=*X�B�%��#�r0�L\�^��p��}��i8���giYz��d�)��N#��qQ��ʵb+}ƕ��UK���;��IIa�SJ�n����_tQ��%��܇�?i��O6 a�c�&{>��ځ�p���׿��)ץڤ¾dO3�ٿ�t��Y6o@�	�֩��e��\������蠸0b ��w����{L���'�͡��Y�з�uptt��h]8�F"Q���Ȍt � 9G)�#�q�;{�><&�&u�1�-g�P���`�Y��Q�-n�NѲ;�J�����
�fWc^��sY�8�E*f閠�0/�,0w4*�n"PN����C�\�[���-�A�oǘ*#�Q���k��y�)޾Ӡ����?��,G^z��I�7�����-,�������Y�9�'es��JÙIg�!7d�{+GM��f���\/�~߾�Z>b-b	�
7�`F+5�V��T�R�M�M���_b��&��Byf�h\�J.�؅F"|�:�����,f���S��g��CU�tk��+���C��M���U��e@b��D�Ȕ��|��?s(u�]���C��T�_��QoXȐ��1���i�t�{��H����$z�)AFM?i\z�b����`����5�w�+qYo`l���5�A3K&����79T���#��()p�nq��\��a�f�n^�
�X�`s6�A��i+�ƥ�G���ݗ�E�dK$:���2�Q٫�r��"b�j�/��@D(�S{�������)�7��eFZP��q`��Wg����I�?�
Sہ��.MҢ��+���ˑA8"ė�y����.��e({������'1��:0���_)�����R�����lI���~�(��u#�V>Qr�R��I�D˄�^1�r4xDЇ��O���&���yy���}Z������|�G�O%���KT�0��l[�R
���` t���I��ug�:<<8&����Xd���Y��b� ��H��X/��"���ޠ��֐�d�KG���A=�_+�y��H8�m*�"D�+<�p��~�~��,����j�H�V8) ��x�����4)�)㕥��i��Bb�`�7�<�O��ly�a� ��P8��}Z%���h�҂^�Q���ݟu�ԕ�:�Ъ`�ILH�x5[���b��S]լֿ�S$�+�ǥ
su�cta� �U�:E�4�N���)����r����=&��՚���r0��JV�O9�������F6"�1�a��X�7_���ۈ24m�5��;Jx��n�#MPI~9�8�o�v(�$cq�=W��	��Xx�y�6�S8�iL@��=:���RC*��'yԂ'̏�*'w5H)e�%p7��G����WL���C�f���e�NH�3B���UL�����7�A���"���q����ݲ����Q"OC��l��'@�;��6��H��y^�J�O9��5�h�D��l~��{ Ũ�]�A�;׏0�i������J�Ft�4 -&9Z�D9���C��R��⟛��%�l���uUq�q�I��:�O�!-�Na�R�0@�kx���A��l��%f�-B�(ku�8�t�8�_^�P3���~+u��
&���b���cB^�)qU�,���$*2?���rn�*����F���2eU/��G(��c+�xJ�Y=�?����'�&��$V�\yL���]Sى;�8�?� �K���I���;�G��������$�G�M���MVʲ��@\_�[�����(���4��P�%�,B���KN��R�^e��L���n�����a��g�H)O똇�H�K1w=�<�*�����a���;m����L}.0�ﴐ���.�,�
��{�Àn���X���i8 @61�atZ���\�0ڤTa:�'pw4T3&�Y���!Zr���M&%m
��nR5�",U7����㿫$ep���6W��ρ]Q�2iNfWB� ��;��Yד�V�"�E�9Xj�n�o���x�e�+���K��gb�`$�겂�s8h��q>2�T[�o`dʖ�����k��Va\�[5�s��pL�?�3�@6���W6�C۸:4��_��}��?�D���\ )B��8�v�*�S�NW�Y%�k���V�]�K���>K^�>%�@X�3�K+�(��Ŋ���Z0����p���q?A��S3�~gn� ��0����B��i�[%�ƈ��?Y�-�LIG+,�br>$<�k$1H3SR4����J�p��uywqv�O�U���}ְǚ3Ι*���0j}��OZ��(���Y���S%�k�p�r��k��
��_��ֆ`��s�Ć��"�6'�C�r����
{k!��ȦeaE]9fY�Zl���O�cKp��=Ŝ�*8�� 3��g����T�`c�ݦ8����*�H�E�P����`�a���|,�JT�U��o���N�La*9�r�Ħ<[�y���<�o��SKTҹ_�b ,+*�Zl�����E̾7ޱ��^9�)>��"	9@��[;��CG<lձ'��]9�XZֲ���)�R��)���N�J��"�f�����f�0�wC=��q�gș�W|k�p�m
ROO�Щq�I�ۛ� ���w$�9�b{qo�z�gQ���\6ۢۓ�@R	r9�43�2����F��l	Z��k8@�0G����I�F����䃨29�z���G�!C�'���	)��)��L�щwRz�:���w��H9xu;=�T���`]&c�o�K�|:��yF��Ē6�8ޮ�%ˁF����E�\�'.-b��lؒf��X49���t�L�0�ʣ�B�|r��F|�)=�ErT�n���@Wo+"$�i_�A��Vx9��f���ݘ�޾�N/�$	� 3�9"�4Ǳo��]���>=��au��k$�E�-
C��?"��]þ���"ׄ�<�ؽ�r�b?ƵT��x��wF��n������;\[��;���lqBq��~?*@I�X�����ܪ��1�,6�l�k����r<��n�Y�\5�: �l�0���(��_TG�g3�v�kuh���z�RCW����oxC�����u�����#��/k6��� ��>�	<j�*�Eu\c5<�Ø����m>�ۼ���f��4�zAĚ��?J�����0��{v�0��diG���I�|�^�d�$�<��|zc�(����d�9��&>�]P�����Mļ��v�IgFᨯ���6)%��d]k�Qk��p5�OM���i���l&�ZA$o�be��b�	�J��`۩�>}�7���X� ��0=�������S��i���yk严WXYr�>[��v&��ʚ�?��Q���R�~� oɞ�4��S�m9��Dsҩ�D�i�F�4f�!)܊��Žgn��x�z.��$�{�Z�~�n�W���7�3��3'��l�j��>��+<���`A� +PB3�� "�j)����*UZ��p��s��儡��!����mx�c:�v
z��"=Nk��Q=��O}�����>nT�)�L��2��2���^���۶пqZ���bd��0�%��+4�r�ٽ�{#�zyy�j����J8�A���/^����\
r�T�8�{�\�y��I��9�&�EW�a�ŭ��	n\�X�\ަyI�v�%���M��m9jV��52�F��,���y��秚��<24Y'�M ̋b��#�ی�h�#*N��ˆcA��~��Mv��=�+��%;�6(�c�u�S}ѱ�h[=q���#����`h�۲�KJ'(� ����蛽��"]i�'�R��_�]��G�5���fµA��h��p"����܄�[��\�Wu;��@P;�򦅘+�9�K��rI����UsYi�$�Y|��} <d��8���~�M3��u�~ݡ˒�²�ѕY��I���_j b3�p$��P�qb���� D\`d�L��� ��d^���+Ó��.A,��4�B��!D��A�w���� ��j�E~�S�$��T���֊Ԥ��6h���j��0�l��
�4Yh�#λ�X��(��w�,�v�X4���Kט�����&���.G�<J�m'q�(9(�/�a� ���A�ǳ�����Z&^�k���N��h���>�vՐ�����[AT�U����M�8��'��׼T���H�/z�v������q���}� H�&�/y���,ORIL�j�]l���c�2l����k�<��U�Wɦr�P�DI�I���e�qF����߈u�4z
$�of��ZPm�S�t��>X�0LC�ի�֤;�Rd���GV��bKN�XE�^Lt߆���DӴ��h��<⩪��}/ŏ�Jnr��F|�kk0��^�P��U�ʝ/�
2�yQ#�E�M�A=+r�e��D�����`c�MON���s�Z�ƹڂ�(�?=�QI���^_ru�6=<����*�J)�(Kܼ�#B���\V*WDo�aJDp�a�_��6^g{T� $�&���[�?�Y��f3��; �D���)���p�z�kK��d�AE��@���\��d(���Ϊb�'����c��G����ᑤ����k7�����X��W�\NVѸ$��-o7s幩>�ؖ*_�\��g,�|yx�T8��V�PY�u^�T�W5Hfm���BEWg�Ҡm�f���=j�f4|��0��� P�P�.�bY'��)f�&�i�HH�o���ݫ�UD��{\��"N�l0�\(	�7e����ТF�$*��i��m�`��'�F7�2���
#�:�t)M3�ɹ,a.8b��ǋl	�q�Y��>K.g� �����^��������F������x�4A }ǟ-`�J�x:xUǁn ���͖ބ�s�O��{�J�M���zS��ܹ0pB��]q�J�Nu�ㅔ@{}�"D���8�����mB7��?�����rr>���1����-�`M+�B�-���v���2��OǓ�؛� �䑲V#}�%�� �"���D���7ϟ^3Kzg�P��Ԙi;�+v?�6�x��|)E&L����*	U��������鲜Jso(��f�$
�30�m�/|�hJ7Y�|N #�H@=��B!zIE�����	����N����D��ZG�+�G�^��D��T�p��K,�i|����<s�w�}ٓ` "�.����O-M�\
<f��G��4vȕZ��fC���-l�C;!�
4kV�a�}5?t�P���3b]��ؠGR��k�o,rc�#��?���W�I��HE=���u�ѩ��[Y@�����^h�k'C�%�A����HE�4坝�_a��^�b�2/�0�
cc�%71�1^���1,�@wC��"�M�%��oáܖ�VQ5HtuPcB��ҝa\����\�EoI\]=��`Mz}�"X��D��Ri��tB�?�>���}�
���1�1�N�+�f��qK�<kgT/�L�So^~e���̠2���̴tP��zZ�i����/�G�Y��:f��#@r���ʊvn���+=��B��̉Ϧ��<�����h2+��X�	!T]՗��2���[�y+�u����������[���U�����T�5���v�ތ��_��[C-TJʬ:Z�y�Q|��?]�[!��e�
���4��N!���0�Ds2���S�B�)�*۶ {��rgL��U�U~wK��R?��d�*��}dK��)q�C%4}�L�-aY��L�nJX�kA�p�5����n��  4��Kǳ쟥�p���an�DL�D�������ߒ�:iTk
f��7����6N_�a}G���C�;{���Iz7()�)�}����<=��ז���6yNJr3-3bN�Y
���NtYϙ���9vivq�odw�ډ{���&��,��ַ"q�s֤�Z�n�Xt��h`�����K�V�I��2���Q��C9|�e]9�m:������φm_ܮ-˜dE� Ĩ��|�����=��҆!�.t����x@z}߽��`�.b��!���<et�m�d����M���oS�d��p�3��2�<h%�)�!����W�#�M��f��xTW�;	��w�����]��&������/�KŬ�b3�C}�C��y��e~�	03r,/`в�����V*��ZQ��o�\�����W��+P T�۶�]u�M����f����}��[@�i"��+�8��b����9��ey�x?)>�`��+�]J������[ZS��R�B%��HOy��w5+��B�n�̫Gϧ;�~X9�!�X�P*ɡp%���V ����]���xI76*BGT;.XU�@��f��O�����+Ez<�.�r��2C�/A�Ih�O��|oUltN��.�S}�%��%���[`)��`��E�=�>d��m3f�]���	6p�3~+a34�r��0WB���H��LMVɡ�m
7��Z��:I00:-xh]=7򸠒:Ȑ�,3���Ie�}$m_��V��L]�O&S�u��neҪ���֠�@B#[��Y:df���ȇwW�����z��ӳ;	�Ճ:�%҃���}�h��!Bq��K�u��>A��n��h�Qs��@�X��@,Y�����~^�����a��]��v�X�0=eR�k�;�q�]�4pZ ����x�%s��_��7T��Ki^�)�	�a�V�3��t �w1tT�U��|��m���!cR��x�6�%����c�W����TL��3��0fOu�C�pUU�j�mh	�+�¥yX/�\�b-����S���.�E���ʛǇ����{���`�@�������l��RY�^�5�X^�N�PF	����9��[�f�N�`��Paw��� �s��
9��)U�\1�N�T�s��<-F��+E�4�mZD��,�-MN<)��;-s��K0MBb\m�qz��qo�wU�6`������_�I�	n���-E���1��b�Ap_ّݳ��kvF��(��S(,w=%�%��Q����d~�_��G�~�Mv/$ڊ�[�@���V�Ӛ�p�Q���M���:�{��qTD����,��]I�����b���j�C����:x�$F����ʆ���,FEV����p[1�LԾ�\� 2^���+x��w4`ߵf���k��+�u�+��km�ֽ�X)j�����:��A�F>³\#6G��3��J-����	K?d���`L$ʘ��dF��qd-R.���ƬB��*-a_��Yƃo�L�l�X�v1\��g1s�.�m�?�g~-OC�a�v+;����Ļ��������4{���Y��ͧ͵�t�[�+/�5��*��i�`n�&���g��U���\�K�����%hn;��]�|��� �gJJ��ރ4��C OFKE�����zK�������3�����m��s�U���P�B&3�Y�1�W/f�ҫ���u'C:ۖAȪ�O�]I~�8X����
�DzX89��,��
�����	�)�9�>?^y����K#"njtʃ��;e¾���T�ʪ���4��xE�V�ܦl$�'șϪN��[�>/��6�ggڗ�
�E܉��얁��Ԫ�z6�7Fc�� �r��Dl�ɠ.��N�A�ْ��:J�ަzU1IRR�Q�Ś�G�@D���) ���K-�KEE�u�@B�ľË:Z�~.W��.���NHP���$9���i�W��j��)�8����C9����<�{�ڼz�9J�C�Ex�)�3$�q�����+5"�1Z�z%B1;����H|����?�
��&k[��)i]_d��w0�����
4���q���K�����;�ɏ�%N&��6s��B(0?gD�����* E���<�ߠG.�c�eUW�b
:��]���U�%���0��P|������!�΀�u�hA�Pu� �!�U�BLkk7Vg�Zb�;����R`�/|�����i����F���xomNi��ɞ���Ǐ��=��0�ܺ]���j�[��x ���21y7Z�ov�^sk!G�U/l,/�w։�8D���#m7,�+Fa�
x�q�c��m�b1?@��*��>����хxi��km��0I
8�mt�ſ�F?�n2�܀
��w-�u��$�$�L>�
��4+�Ϝ"�����N(�{\�0E�Q�N��A\y�jE����q��& <ÿ�$[����}̖����+*~�����U��~�d���?r�=�����0c9�Y�3!2��>�=?+��Q�!dУ<{Z�� 9K!�����[���#,��Q��Ů@9h�	<;x��m-�+`ȕ�屣�GT��3ome�8��W��K�p�b8��Фi?��� ����~֬���to+ק��5���C/ꒈkR����#D��}��9���B/����>��>P���[�PӮ��Z�=4Z$�R�#���s.���,�,ţ|_X�ǵ%BtZn��.�=�"�� �$��u�zrF<z����>����~a�ο{p�����%l�w 2cT���s�=�Y�ԭp�j�J�f.]�#mI��Je���gL.� "��I0��T�.G�fkg!u7�Ce���^9|�>de$�>���8�����G�l������q�L�h�=�,���m�3M#��2�����u��/V�I2Ʌ����)Z��p%o\�G�;�@5_d�+��m��\��oǗ^�8��8�&Q�iR��;ɸ)�}�r8�V���,��/eC�5ӌ��p���dR3�Ù��k�y�p"Ӥ�K?;
l�EL�Ƽ� �Ť�G��P������L��|]�}lb_ǮZ�-���S^��f����W�<���{ϰ�wd���f/_�Ћ܌u�<[�H�F�<#M�("����_�J%'���I"�f�y�$�����]�Bç��˞�\H��e�о��'52�'\���|��ȓ6^${����@�%9X?�.Nh��n��-�O�>�)_�8Ќ��J- _v�}���ub�����}��c��W����,_^(+��7Wc�q��S֥���"6�p=��S�
qZ#!��Ǚ�k�Ң0�u����g(�W��a���	�d��RӤ߳$���$vw^���Mz0�.��y����k�Jl�m�g$�4ib��A�vOt.��N}M�лٝa9�_�xl�;��6��������%Ƚ�r�:�D�'4b���)ɗeMS��t�ꩵ�]�C�%�3���b..����0K� �'�e�J\�|��D�6o[�3�A2:��0��	��'�t��m��� @��Z�yY������|���iٛ�bO1�k\��ނ�o�:x#��<�'a�w��^ [��7�jt��5����U���hH��e`t4�Q��301� ��Y_J�>���[����e�����ӰJ*$AG���&霚 �Z�^�Sx́p[�B�Tr�Ӱ4���f�y{b��OՀ���b����=y0�|�����e߯ ���%��2�N�e�z��$6��7��=�C���y�9��K	�7��V��UR���\u��:+����2���>� =w#h��f�6�A���
��nC��F=�,B'���RW��r1�M�P�׈h5{�:���4� )��0?WLȝ�Z����h3H��Kk�Xn�O�Ne:��$6���Ҩ�����Ҕ��6��P,��x�Hu<�(D*��� 8�1�9z��.3huk%Z���\��k�
��Xk���5��6J�Dg,�b��A�W�A��b%\x���1�3�W�2�J�q!�Q�q�	�R��K�,���'@>Iu�����̳:�9fM�޻X�z�\k���+b��e��V/n׫3�v�_�|PÌߒ�6Y+A�G�P�T~�J�-@�FU8�t��=�nl�^#��j�m�gf��P�D���ѹϺ��uv�o�W�ˍ�l�IQF����S�/��]�b�CP\�����"���	�Lf��ߓl�s���0�{x,��kn�ٚ�(��ntƳ�58��6��@��;-��g3x$�#I4㑄V�x���[cA�1AL8q���v�Ш��y;�Y�#�T�}Q�&�[�`���>��+η1�߬����c��:�މ[1�<����Y?ǎ�g��'��ߺ���g��("`1a��Hj��s�7�3h���@6��j	ץ5g5x{'����c6��N�7��-5��$��ID�"��ÏòZl���ڈ�� ����3��K�@hd4G�ҁ��
���W^	��B˿�g����O��1����D�d%�5��.&�-'恜Wx�S	���t�z��o����K} ��a-^R�o� ��b >�f$"Tc�kDywi���qW���1���đ.Tދ��y+KUD_+�&t�x`|��V����_?sQ1c��U!~��:!���cD���Y^y5������Hel3�/��2u�}l�\d��@�'I��P>��l�+��0r��"�-�DA�8K�-Zd�@=��oWaז�}k������)K�t` ����a��) _� tF�k:	�����\y���"��q�"���5[�r�eւ���(�/�u�We����%`t�[hs��I�����W-U�EO�ѯưkHĂ!�h�q��~b�K�Y�>���	��tD3ן�ˑ�L;a羌;�>�/���D���/�����A���t���*�I�Y�H!�^�7��x�_�Z,A��sug���y�d��3GJ���^(}����5;,�6��SHsFYF����] �g�%6K=Ud�c��!�>�<�����lH�o�&�{����`8���+,��p�t�=��G��w��r>#Q� t��xѵ0e_<�y�����
f�[-W�0�9�w@�7k7����ԪkW�ln,��,�Ȩ�7��CRuB�^Y�DzD��āss�����sn��}����|_� o�!��.��sJ� X 6�ü'�0 N0��Q#a����N���g�J��9B���#ǥ+s�&ݤ�E��Z�O�[�d���7���RU�X�\�B<��O�-���z���`>D[n������|���:�}�cM���\=oF�v��+9�ɲ��ײZ�_8��jZ�)Օ҇(����2�U���à�1��p�.�Tŝ�/p�W��I��6�q�8�_�d�4!���������,�m����̶8; L�%���@*�c�-�����~�n$�p�S��i���r>��ZT�}��T��#.f��ڱ�;�p]���B���XQ�f��]����@�%��r�-G;��l���Y)U���5�Г.wM��ww+Ie��(��s{��˹�����j
- �F��,U&m�w�7�D��,�?7���?��S���i���yD�f�����u��������K��P��a��c���ص��Mf�\ï��A��i�a�W�}Π� ��gu���[���2f�����G�\J<˹����]�/Tv$`����$d�C�������pz �9j]׬���Q����|#�z2n]��c�^2A愙�I���K3��`5�tgW�1rˑ
����rM�����ݠ�u���?bv`�� O��p&Ԙ��D^߉�i�ħ���j/d��
l����g��k����E��5A��u���)����Qro����9=�~�|pX�R�8e9d}�v��Fn���o�����5�C���jk���	�,B��c#3�,sؼ���
�ƞ]j,���g䂄�\h�O���b��ܜ-�y��~5{�J:��V�#���Xé�h��C�碌��c������b�%K���J�w�j�k�����"��:4����zEC�J�TI��"��/-�,�u�����h?]| ��Z����N��c>�QC�B>���J��@��,a�o��C��h�ؓ��q�{��H�����Qr���<(�m^���Q���&���@"�|�*|y�M ���3�
���쯕z.�S���IL��;R7��M�l_�藝į�B�>�X�=X��lG���L+�����\��WV� ��D�2�1�_�I0��K��	�3�D�V)�Ҡ�~�WOq��bM��ES!�g�v0->�nb�3��ț���'��K4{���>��u �Qk��� k4���+���j��+@PN�?��Ӓ�l�B"�������U~%����n�PB��vy� �:��������rQ"I���kx�C��#���I�ݟ���'��}�F�+#� �Sy=�Lå��{����g^Yo*�|�n�:yЛm	�	�y�.#�v�\2�W�yZƲ���n�v0����UW�mM�X��������F�ڻ%���[��=�����,��Zh�C�;)h=��u�i�,��ʹ�h��:���#S�:R���{'�۳5����ג�f6e�]�r�p�l^S@�xUB�X�����ݥ��|=�_�^t��u8����4��9j����}h;�ξ������"�zi�	��Ɨ����	����Z�?|�%Yz�����Q�D��Kƞ�1p�T>�F��%���{�j��QN�b�	WJ�<�����>�z�/�����w�B�¹އ�e�h�z�G;����a�H�'̇fL��e�+�ؗ&�5<�v��!��Zwד�	>�d6�M�=yP��g���?�V���hyT����`��<�c�9�n,�3R6^/�L4j��6��KG�-��$IpսJ.���K�0B�^VKꄇ�W �%����e�n��qa��fr�d;�C���0��'�~E���Rf���w9M�VV�'�?f�%��Y[�m�?r؄?`�F�?�?�b��`F;p{<�]]Ԩ�)��r�uN�2�����i��%���U����Ƒ�1B���c:�4<�0�r�w�,m�{o���@��B�~~|ԍ�iօ�h��n��2������A�"4L�ᢨ��T�&��_�2q�,'͜}�}�nG{���L�I�� ۣ~c�l0�1(]����a�Őqk��K��T񢅙?Z��0w����9��><��CȞL�3�s�:���]2�>����b���3)^x�|ƥFj6��E އ����ӎy�W%<���V�C �w��
�֋e���4z�8�n����mp�߂�r?�e��\�]F045d�O��{�N,�,o���!,p��GAa���j84e��W��!�KE[�ݠă�堑k19$<s�KMm2�T`�w�֕�L���״��5W��JG��ou_��'�cTR]��b�*��1V+��	�H��>�c��8<�=�X�-�K�LtȦp*�My�5&poT����i,����0���x*�����_ɅM&�n�c�c�}��NK�� wΘ���z���}�rv�?R����� �I�&8��C�^C,4���X�	Z���}- �ư�g+�2����e��#���M'[G�k����!�w2ܿD�Y�c�5�/��kv���x�
=={#	�!������d�Ϫڍ�Bj�;� �8����Cz�p�S�\s(ē>���� ����Ð~p���@���u���=m�壆�ӪT5,6�+]�#}�ơ�������]��kTM����'��k�O�����;���|��6|	j��f��+d{��K'7&�{޺p���D�n�.Z��CҮqj�����G)~=�i*}y]Z^��2�V�9u@0td�j���hm��gܫ�qVRK���~{�P������3����H�TJ�-�m��c/�{��Rޅ��F��r�<[�T���ÀSa�wM�"@<4dEv~6z�ƌο��o�K)LE,NFV�>Վ&Qv���p��O�~� �R"ͩߛ�eo�sj^;�wG@���?W����ՙ�j��Ҹ����MD+�	$�S�5�H(�{O�H:����kn8�R�l�_�-3v��+"�R�-bӣ��Rr�mE!� ?������(:��Y�}��U��F���. �KQ��\T5��jrQ���,�� ��t#���w�Y�����;X��M�	o���xX�z2P¨#�R�`�*Di�x.h�J�[��i�O�0�ӝ84�@9�~dt�|�8� -�́���D�Pz�v�H�vPy��xQ����s'���ӳc����)�L��E��N5�5��դN>_�ےp�Kܾ|׶N���D�&�X���/8�ebL$����	
|����6y�ס�.�KHa��u��=b��O)���JE0K�U�_��u(A�)�튎�R��b�H~�[Y�{�4R�*��q풑��O��E=&1֮AI6��p��!�����$�f�'xct���G��<�rƞ��K�	�� ��k������{�Zw���+��ʉ`d��CiڵMK]�V�R\�zW�S������� A��ͬ��HI�k����b��>G�A���%��փ���OL��I�1�#XG2�{������-"����S��k	���o z�}8ٲe�P�	۝(?��1��2.Q��
�[9�zڝHm�J��*h7�u	x����c_I*�[@s�f@q�}㨛��c�A	0���{S*��m��Y��T*���i����'���g���H��j�@��3�95�7�n�{O9 �N	�(j���7��;��	yv��G?�{k1�b
����mI��4�_�L�8_�Bg���!�{}ʸ+�]�x�}{w(�~�fg��DOnp������A�B[��7���:؛g���M�R��&'}t4��O(��i���l�ʻ������i�����4�A�1�ʨ�匒fD%�6J+�}��T��& �TlݓHE�r�bs	��$�y�(�g���]E(�'��v6�-'�H1|�[�m�	9��q���첗��7>r����c�=|����V��n��v��+�a�ѷ�N�JK�\��G:p"�Jh7��?�_�}�v�q�0��'Ŋ��q_�ڏ9n�(��ɏ
>R�8�u,�.Wn���rȕ�51|�M�CY����� X�3΍����n�9���#�[���L�k��AV��="n�����䐄��.�C��׻�-�e���ƭ��7#�� ��2�o�+*�7���� TT�b�;�u{�< �&��sL/�N�
��k�M@�x+S$vc��ע!+�η�aX�{֫츊I�x�ȋ����"���vT��U�7g���(!�L�b��ӭ$,�l��8/�*��vC$�f���M����<��*x����<3��sa�d$^�Pb��y�������i�����36�XR�����[=v�t�
�����v��"ҝNr�l�mz�����^$"ݔ
ɴA����ׄЂ����;$���"�˯�����C����>���Ƙ�^~�J!�:xb�{��W�2�ƨ ��x�P;���8�;9���x��JCu>O�JI����C&����_���a�z�F2�E�(=��N#Hw_�ǂ���6�?�sd�zH�*<kǆ���Y��g��2Z��(��).^BL �����R.�x���O������%UjH����M�N���k�,}���"�*�Ae��W�����I��k�3�����d�@�C	��fh�4�Ӿ���eU�.1X���["!1xLX]��s������ Rb��K� �O&�p����h�6e�r��2h��C"��� i�������H,r����f?j�R#-�fஎ@��wT�+z$�3o�Y�=�����4d�ɡaZ�f�Ǣܒ%�4o�&��gH�/G~��ow��7����=�D�\��ϒgbW��w�:������Et=	DoW:��W���jFa�q��ZB�T����tyT��>;qS���_�:B�^mI����.��iMq�+�?�!��p��ޖ+�kR��WL��O��xa�z�m�_���<|&�b�m7z9\^��S\Wlo����˒*6XXg	�2m9��v���*Y�Eg�$'�x�;œs��M�xljp%ǚ�.�֤x��{��_"��DR��u�:0D�y6D���&Ԋ����I`�B9Ō����h���W�%e�����]�|N]Y�w�N�]~�����k�p0��П�����6�]�M��"� �����Ƴ�J��̲^�6%�e搀�Q����0�>0�Z�J�[>�oԛ�F8�7�̤���������dH��7�m��l���o�� @�
3�R�=�4�Ҭj��hﴵX>?��X�xԍ���z����k��FT���q�/5�����Pf����t|��3�Y��ī(��d��,�A�����&t'��9���O&jҏ�ѩ@h��.���h�����g��z�m��f�`(��)�+�<�xգ{�D��Y�>�d�L�k�o���m�Z``�Ş��" x(���J���2�+=r���j��%��)޵�� �}6dɢ�>�F�=fe�alkP;�/��c}�q�0�I�koЎ[H�=��$�4��I��@ձ�9O���
�t��U?�I���X�Qt��CUĝv-�/�[���=#�a��I]u��AboN��x cZ�_�[��R����׋��0*4@���>�qVK�Q1���xo�s���㩂���9ۿ�Ì%��
�k!�%�"~0��������Tp�(7'm��Ę�g�Q"�6���� H8�ᘢxJ����<�*<��yа��f(�)$tz�������yt$t���,A
J�í����4�5\�r�׷��@�h�m'�A�a�/ �Z2v7r��gk���U#H��7����Iއ����+��R��CR����,Ym�r� ���ݞ�D��V����:��O^>q֞SYT�q9zUQ��'����1���U[���8�O�R���v��R��3P^��p��w
ە:�z�L,U�fe��q��P;G9�K{�<�Z'����Z�z$N��=*�K÷���������h��gP��j�w`�1->Fl�����-��z��'z��|?�J�'t:h�~�؄b %����v7 T�6lj��$������ҕ���:k�tS�+K����l4-�)0����r?�G�����"w�������K�Y��+��g��_�Z����2X�	0��Y
(��1�-O��ó	��3Y&8\VQ7c��0d�i�_��֕�wb����i*�w��rE�����t~�hyy<�$��=OOa]0ŝe�K?�c\*�O�)��e�~{��>���ð�N��	Cm  ����;�3�dpY"1��'���(�wb&�7&2E��Jp%u�.�yD�����vt�j�g�!�B�v�3h�x8>Ƌ1bѲ�R�)�|�I��b���[�R>��@��|.��� �D|��+�w7���MZ yXD����{���^�o&������@����A��2�&P�6K�o�rv���F�s?�1#�ƣ�2
K?=x:pJ"ѐџl�-��쏖�`Ek����A�d�wO?����8�����oy��غ��*���Z��jѪ���,��#��{"l�D��E�JD�M�1�����|�DȊ������ٻo��:cj3��2����
�?��kF$� ���L�MA'�t�S��ԐTȜ�cx��
�OCu���8,��-� ��c�r�?阪�-�t�}�ȈU~m/�y�8�s� �����NX�m.�f��
����a��q���b)@4��Ϗ���	��' ���3��d|t���I;��T����y�YߞLTcA���,p��M���ʀ�l�6��\�`'�.�,??�����{.$ �!�Ȅ�y��Gف{��^��x��H*km[hS����W�<)C�]� R�hW�mbw������F���@^�ڗ�ج���ά�!%����I�DÈ�B�2L�.ߴ>�j.#��y��ް��ּNa�#�C᣷(?�G��Ja/�3A��Jf����׭Z�m&G� @b�(���mWv�#��t���<?�\��Y���$*�%�s8��2{+�m����lص���%��k���;���z(O�,Q��8�4W@�;�ƴ�7y�G��d��0�.��b�z��D�m��4+�Q��v]����T��`A�H|��q ��n�z-�E'��#�)�P{#<&�=n�7��4y��$�V���2?�+d��/hGi2�+d����7��ϻ�d���z�����T`�\��t����c{��W����BdJ���֯��\l�:���d�R��h?P�l�
��s�b+j�i���2]�x�Z�\���o!JE"3�G���j6���T�fp�fZw \�I2���[�6������*#����	==B_�G L�ՑE}DE�,�i��t�7�%��o�)9�D�7s�&�	$,j_¶HH�tه�O�6�f��2������y�hFf��� @XxwD��
����F��w�wn|��^�|1`7 ;��L�����=O&����~T���<�
��xm4��|r�Q��!�
,;��&5I��|*a��|v����$�l�t��<E�م�{�I�ފ�y~��:<��^F�i�7�ϋ��U�Ƞv�{t�O����O`���L�嘫�3����g�;��%Ʃ����%�������<����"襵[[����xTk�*n�
��e����	=W�����!��,7��&n[�%�h$�rJ�H[��W�q�n~1�C�o���5�uP�yvWg�o�v�l����Y��("�Z��&�\#�UT�"6_���źf�>��0��l/�-�.f5Bh�m$(���+T�V����b�u${W���2u�V$)�X��bDcp-__�5�z�@���@�!�̌5*���%���bT-�R����b n%����) ������o�ǴLL�{)�>*Ѩ�����3&��Z��/#=h,�E
��̧F��}Į>I|r�g�Ә �i�&z[��e��$�ԋ��J��{�a�g2�M�> ��P�d��a��U��z5w	���9M7���ԍT�|�b��d�kL��<���x{��&�Բ�Է�+�؎�h�J�AW�>��4г|����/Q� �F[$�7�bc{E:�3z��T�cj:(�ĥ�"��%�x�?P�ao�N�PUyI�B��28�΄ˀ^���߇	�C#�,�Á����e�O�%�`"�_�;8�� �~Ckv��l�k���N�Ŋ�1矣��]�r}X�C��%u�[*��l�,�:z�/x�i�8�h눨5I4�L �F Y�\����𭧤eT3�j���ð]�2-ًYl�9"�z �Qs�[K�O���aA�_�'Z7�H%a�6���:��2r��l�����1�-�S�A�*̰�u�}��SG�a&$'�C|E���}�^�Rco΄��P�`����*�I9�Z�{���2��!�-�}���+��㠱���{��0����p�­�8�Q�+N���qu]O'�e��f%M�ۈ�F�D����bZEf�窢l�����Ge�.["X,U�C9����xpf$h���,\�"�pG�(H(�p��+_��.�c�����L�B�5_�̞;� `�#�N��H��%?vA#�ž�;t�V#F �)�)zxf0f2�T"b/���F=�q.*t�	y�v�t�GƁ%��}f�0�
�Ѧ�C�n^��	��Ut]�;4lRZ���s!6Wf�3RL�ϘYU�&�I,�h�7v������ꐠ����S����vJ.���v���A�����K�$�g=>3����E��Q��!\��:JEb��s���P���E�:��xA��������:�T�Zi��OeCW�7��_ϱ�c�_!��T!q﷗�v/�UtHb�1_zv��"�b��V��]��X�$.���Z�Q�ś�l!��p��g������-���9J]șlQ��k=Щd�Z�����դ��gv��z��^iⱆ�ع�{"���1�u�w0�=���)P�Ӗ�y���|�|�g��k�������	����i�^{4#�m� !�q�Ax�g��-�Zj�4�� ����QV�#���k��s�J/��n��)X��b:��e��|��hsOZ(���>@G��[熹C�5A�����mގ(3��{ȠOl��qdr�]���t-�Hon7ì��eg��Sf?H��JFVBg�|f|�g��Z�ɉ���0�S8ݵ�+�N�p�C�}(�6�ۭ�y0F�v,����d�㥢�b�4e��\�P���2�\�أ���@�_AI���R�Wϐ~j&�p!,[LC�E��v��Гu!���m�,W/�,.�Pb/�,!�Fͳ���ͨW/�����s��@�O,�yy�T��ޱ*~��5�r8��|���<��	#��%��h�$a!�Ea����&�}�b:��'���F���{�"�����T�A���h��1����t�*��n�Dub�ݭ�s��_T�Y]�c�����$t>���e	�3 �(��Nw�f��>�A�ᠸ��\@����3p������H��[���پT�@�p"}�K-%�!��<�(��0�Kh��LK({��L�<������m!��m�>}�ҠYF`�������4�
��i���泽7	�J,�������Y
�u&���T�&"�N��s��Ocu2�d�YT�ĶE6�W�W	�;���_H��&|`�?���,�4BJJT��?�U"�G��7���b��ej�'S{` �ɲ�ET��;�k�:������x����,�w^��>��%�N�#���������$T+.�Ub x�p���VF@� W�1��Z��L�@����f�~�a�:6v3�i;%S��!�Ğ�R��J�L�-��?]��N�t$������F�)#<��1ܡ�������G�����E�["v�f՗9�����J�cYsV^{�.ܧ�1_�㩥�yaӐ9d���g��u�]���xp�{����PD	��㜾�r�Ӱ��>��Y�eУ,	�`�7U����?S�̔Il�?���N,9xn��������UmO��/�!�(1�����|t0>~�$)�,nZ|���W���F3�A˴1�nj�_���_�B�W/�ڇ���T}¯��W��	N��,6��~R�+ኾ������1�B��̌��:L>��42��Ľ�}�ABS�Pǂɟ��w�����	Ap|��`�w������P#�S�=o�8]���&5/�e;��,�=�YZ	�Ciul��������`�eA�_����֩�O̅)Ytm��?P�}]WD�k{1l~���,�ЕZ�f(q�g��>F,�5�7#KW����� �V�"ax{�J߱��2 �ɾ�M��C}��tj��� p��-��D>�+-UZ��Y�O�F����y<�mk%f��f��6e2�]���Z`�V�R�B����Lf̷��{M�o�'ȊַX�t8"�p��-[0�j���D'ƴ��w��#L�<���]:���J �j3�ꐈ��Y���
��"o�S��_Ņ��ІwF������S~"�A���*�g��܀&M����T�3�X��$N��d�Dp���)4Yǧ�[B�PH�/�p�z���j	�-��sZ�yK�I�FB	AH�pEq�q���u��,z��#	~׮��[H:�!���J�2�v�fb�/|�Y�8WÍʡdr����i�(��0lװ8oU:��e���!&���w��/M��V��w$�0j?�[���<���#�4оx��r��B�;`��_���L�%�@��2C<|� Y�Z�dj٨Q5���+wjSY��� �>���,Ud#Z��i���q�b�'����{=]K����[V��<�qSA���B�u=�5�8�갰2(E|����KK����HP�M-m0��mG�F�+ٓ�	/��(�iΖ-��&YC]<6ˊ��^}��]�/�m�f�û.�B��;�ݒL��|i�o��c���2�qU� �)v���Y��cs�(1�;�x�)CO?�MD_��V�0���s���xCF>�2'���ecS9B��@�ݙ����b.+t�=e�5��\N��&b�H��g��޸(�?'5}��7�\��i�7%���&���O��."ҧ/9�x�@q� ��V!��j�A8�?�QEוs��[`�3wG[���3d�/W�?����ԠR�_���V���3��M��b�g����$�L�` sv���xE�+�'�D��
Q�|Vb�]�w�\�l,~����&�B��Nڧ�Dc��J�$���0�:���[3
0T.L�B�����wC��S��h��-�c�lA����j���=���Y���(��*�,��d6q��{UP��}<a�R�F�<����<8�Kަ��I��_Kc�$ɏE�"d�2*�
�[�ף�nʽ�>�Z!�rg�"��J��lF�\�CH�'�D���:���U��h)�L��Y��{M3�����(�=�H'��)4�hD�KM�$���)`�bkI�)1��.gcZ��n8^����xl |VG� %!��p�Vyr(�� +��U�15�P��r3�꽪]�_w�Š| �5ȿ�H�@�ÄL���)�3�r���Ǆ��Ӫ2��E���3 i̶�싣v�A���I(.�pS�yr8\=P�C������4`n���� ���'�Mف�q|f��� ��!q�A&$G��l�[�ό 1�1X)�?�:�R{`�~'��E�����#`umu˛u%�#���f��t�FV@=�}
~�)lI@���q�4�ާT9��U˻�WN��d�e�絳�ʚ��B �m��Y��?����68�u�Ym��s�Mq{s�4k�lH�!�ME��D��0}��u*���g2&_�y\��I�������>z��Q~6t=!P`ǘ����U��:�f��h�2ǉn��D@���-G�F2_��;�֘��1X4�%����m�\H������(�F�	aVr��_�n�����M%|6�}GQ��0�VtcRآX�ޏR��p��]��W�M߉�;	����(�(_���rz�8����1b�k,qTn1T: ~t:����^��lz9hp�YM7���2��g8qD���@�[�����@A^Z���H��5�sb�j_'N/�.f�8P�y�T�j����N��G3nܡC����E�_*��s�t�|nH�4�-���}�iDoR_��F�G�і�Z��͔������o2�p��IU=�w����
t�Day�p�V�{��OF�OAU�����h�1_$0b2�����=fYg��\pN�W�B�IL�O�R]������v�={���ןW�S�Ū$#E����
?�N��rz]��ȧ�=�ܯ2�ua 2<�9����W����p�Ŕ�S��ɹ5X~V��Eu��bg�Ъ�k�զ���Ұ��yůӽ�\��YHe�Ri���t�7�Y��L���/���-�dpM���i����(����4q�t�[�Q&�0BB�td�sp>?��U��8P��P>����%<a�kP�s� lw�$�itp���e1���D��!�c�TE,h���Ny���n����Nē b_��~vFM^�>_3��kCx�=��5o�mtF�i4�����b*k;la|a���P�dy|�Rt����4�O.��j�����Ce
�vn�;�a~�?~�#Mٵ���<o]��� �~N���󢈔>I��f {���m\����gH���������qP�ﺫ�}Zb��l��L�HSݯ�y��<���׶JF`Z���`����z	=$|G%��	�$-.̩v���q�����ډ59h}�e�D.�����	ȊZ�Xh&�D=��v.Q��/���g�7�����v2X	9V�#xy�����0z�I��h�x�߷�8/ǂu/C����"^���/P'�c��3���@�t��*��Ұ\����@Ս��B�U����\��d-f��!,Us�n�P�ӝ�&=�V75~ŃsD��tD�(�O�F��N����K�E�;>vF�̶�jI��9�p��I!lR7Fz�g!z�t�^Oq�Z��=�wD7���D�u�,��h����Eo����ϧ���:��� c�{�<�L3��͆7��9S�Xiɜ	�YZ�e6T=z��4=s��U�0�x�g���[1e�9U�M_�l�����<z��ԛ��ky����c�rT���\��>�/�PTC_duO:�7J�W=:���7�*�2�3��d�ɘm�^r)Q�1��2ͅ�3���n>A�ѮsoS�x������l�%Zv��."͖H�8rs�;�	/7Y O3[�_������҆O��U���C��-hH�$���%*[��ߢ�/�0J�	��{G.��5�b&�U|d٩�J��h�4�mۺ�v{����L���u�!g�Y��^��a�2[v��H��ȼӖ�,�������L�u����z�"p49E��|܋@�� <�ֽ<S\;8�ò 3ˇ�T��ϋ�fn��;�����ag��\0%�=�/m �0�0bd�D�v���{ܶ�{���"����{��{�.t�G]ɿ�����U��6 !����VG�G�$p�+�N�PO=&@�=��!t���](\�v�1�&&�ߵ�s�.�C��Wg��X�>>>����@* B m!��<�v �q�>Ջ��/]�Y�4R�!�E����Q	kݯ�� ;����轾��,-Ǉb�c�xV�T�Iɕ��L�xo��MG?���Z �vo��U�x��fw��������e3����Ğ� T3A��Ji�����(U0��aXhR$E,��WRC���R>Q
��SǠ�6VV��~�2*��B&���yn~$��l��J�U2�L���Lп͗�@��c�(1m�����^L(���\�A:�i��0��0OxGY��bB@tZi�kn# 韁o����C���1�Y�����i0�`��*^�ec�|��2h>sN�ꊠB��h���	Ck���ð�1�,�r�"s�"h5�~�����m<������DޜH�(ҀF��l�B�;9���pza�)����嫞d>>�duxѸ�}n!EiϮ�����7��Y;Y����x��F�*C��KϋE��$�O,�m|�D�W�@J��և�����8o�h����M&�u)2k�1DU��z@K 7S"�4d����'���V�uZ���O�C팮Aa��Y�m����l��_��Ԛ(�ًC�(�6�WlJ�FV���0���׷{�|����ű��y
��SגR(9���N�t�٬��;ܽM�=�^$����;��Hvs��IW�G���U�3+[�ʧi��	 ��e�����*��C'$����� ��JN`�_Mc6J/uf3e�� �S	z�O/7ȸ*�]djd����x�6޷w�����qo߼��
a��T��F�2�,3�o�PT��-'<�%�Z��|��/�d֮���>�d|����� o��H�sjW�,~;*GM���}6�M�������P]�8�b^�}�D� ��HF��s*Q�[�f�@
�������J���Y���ԓ����kU�Z~�:�R��=i��rg�
c+-My@X3Q�)��#k�E���ښV���;]���{���!L��& �q?�e�k�w0Ď�+�� 01��S�gZ+-��z|q-��)C��1�	|ۙ�s7��$��R2l97���BY5�@�U4� w�����e�:��M�n���ȗ���u���)b�lNQ����3֙W~ �,�J�_L	�mv�U�W��t3TR|l�SOݐc�c��}�A��^~�!��R�L�}T�8w%��y�ύ�r��ʐ�}
�wN�Tmt�VG�w��qf�5bG�\��<T����67k�M�`�������K��L�W]CX��!]�r�Y���q��P.��ι��rN�woA�4\��K�S��+VA|�~,�-Oz�z�.}�D-O�������u`iT�BoS�d� ��$D�m��$M{���*7Pc{�ڿ��E<�\���#8�Iޚ�[���o�����	����fy��b7	� �Uu+>em�{�ɠ���{d���Y��Q�J�p�o@���s�*�n�GS�6�J�=�r.M���vڮ�����l��%F0�Ƽ��~�"�LP\ws$zX�2s�;���G�̍)�/�'�lR^���"�F�����^��z8������E��ҩ�Jf���\t-h�@�}�>>^ S���2j<f4��@� ���4��òݮ�᥁x�@Ĺ�^�3P�V"�-c;�<�d�m�&q	J�Ӹ؉w�Q<G�§52j���퇏�8�-dL>���)��(�]
守���Q.���C�EL�k�k4F�\��V�t����{�����D�ۅ�d�g�;�u1ڵ�ǌ	:��_����2�)^�c��$�����cb���[R�_��6P��(:{=���#�uu_K�m�Vl��jSI/)�r���x��!n�L<�z;�,x{kc�v>a��{�X�r��.��(��ԘM�M�ǝ�D�0���tKA�~��>��vmrQg��l�UP��p��і�9n��*��
��ͭ�\2n�S~�
�ᨒo�b�h��b�X\W���-9�L�� �0ڗ��̃�>.=4i}0z�a�ئ�^9�<*;7 :���5�@��r�KE�fVs#��=8�uy����.��[@
U�H�F�%C ���!�u���t�7@I!���#''�5����Rd���C��	�0��3sz_����Z����Nb���6��ΦY���)��A�Z���+�cJ(u�����չ"��H�h����
ؚԼ��EG����]=k�ϭ�a�v:���5F�����m����A���\�|��,��^��˃l�po��Ȣj�����*�5��n�={W�,|�~uJs�!Gx�NW2�'�L��y(:xax@@ry\�XAY��u�Hf��+��ߚ8�G�9�pV)�E�u]s|���z��E��ǭ��-Ԏ�޽jȼ�cX���^e!���t�u�}��qS|S���ÌC/ٝ�v����x�����&~'����k֋���b��s�xw��'Yl�����{/�	 J4>뙋��'�!���C܀%�� ����2��`>�)�����}�o�d�,� �i�n���ުO�x3��LB-�=^2H2�͆�����H"-� ���A�,�Xm�c��<0���$�BI�	��L��� ��.�ݥ ���I?�L]����e�R��+����Lf��)������x2��Zg
��;˪uA��n#퉂�V�}���p���R���`��0͸���%��7@�E��͗5d-ߩ��=���� �,s\���/o��@�wO��N��H	��q/Ih:[n���!t�����E���8�$�a��V��@Q��ZL�\�N;7�7v_k3-y&CjZ'�̿�p���*��E���2��}#1h��=FxE4d� `��J�\��>X�VJia�E�,�}��<TV=�R�A5Y�U� ǝyƜd��4/�I�����0��n��@
'���;1Qi�h��]�#�o�^q�S�uLy�gQ.NV�֤������l)�F�AH���I,h��-�x?��<
@\u�6H�fN�<�I�������*�)�j ����]Co�g���-�-bq$ @�β v���Ag�2�r��-*I�j�s���n�]����{M
rMe1�O�w�K���_z[���{�?٠�:PF �>	���W?�eσ��ƅ�ט�Xz�3u�"ަ���>�+Nk�C�]���zW;�)��=o�Za0!i�<)Km7� qw&��ʹ�y���1wmC�0�+Hp���f���'�~��7�f+l�I��r?W��"�IGb4��S��-��������q��EցW�ǯT/�12��*�y�1D����Ҷ���s ���J`9����9�;��� Q6]<l�e�L���r@[%�Yt�,7�R�j���_wL��Z�P3�"/
�|̈�{��R�]�����R�V3M\�G	4��=���Tj�5�\o�)�!8�f�7� �����>R�߰�'��T$�e.�al����f#/#b˱�>0�n�o,��t�^�a�<�.w6U�
`&�Yt�F�C|6��<�J
A��[p��CVK/�P��!���)c�sj˩r^-�VYC�j�C=�<�H��e����2*�֨��-���>p��BSbVY��F-���sl���HA5����c=
�ٖ��_}�\P;D8���rn�#ѳ��Hk���C,芁j�;CZ~4nW>5&YD0���*t�4��k���@6!�xB�>�.��@�+��!Z�k\9dC��l�av��A=f��n.�����f�͈� ���dv�M�у`Xyݞ�"䘐F�1�k�,��	A�`xN_�>�*�bj������a�C�9,K��je�āQQ�Ч��e7\LN�L�;n�8�S�Y5���c�1�� �XO��j�R���Fo}	Pvze�>q��sX"�	Y\wɥ�{#{X����[�w"��т�8�D��[F�������8�/�g��tB�O�է��0#�ed�B��ڃ��G�6��b���v
1��Č�\
"^�T�/���	�m��6T7���V#$ˠ�4�N��Nc���`Uࡋ���^�`ӏ]�i�١r���~yȁ��TRƲ �Q�����j��h��2�fm��s�7��{t7M0��~j¥�j�#a��S�,�a�Z�r���ޤt�~.*R��n󍂾t H�a�?��*�N�*qx�KZ �QͶ|�
0�o�=�L′�K�!�V�½�v�5�X��&��K1�f��P9<�B�V����'1�d���=��]@�:�%=*�+�.�d�
����[��DS��hLϺ��2���0�A�n	�4fඖ#z/�T����mږ�ʈ�pG��ZZ��g��#؞����Ovt��aE�k6Or�Z�� ��y��&f@ۈ�q��̗�T�S`_S|�}=�F����4}2E�:O��̮��jg��>^�v��FN٭BuS,�#痷�:.��1��2�[R5��\|g�L����%-����ک+��2�@��޿� ���>��w}�Z���e]B�A�����[�x'6j�eɀ���9]�&�ץ\O�Ȍ��	<p[�2��P�
ٟ��K���y��K�&����5�;��B"���JJ�F�:�XO,���S�i�8�P�?�z/L!i������)WL��_�R8$�<9�>k�%��&n�c>�V�4�m	wq[�W_�pZ�_��=i�6�s�Y�8�.�䃼��I��q�֭��%n'�!����;�>�P� �f�Τ� �F�8q&�]ܚ@�cXa�4�K��1&pӧL���)�8��4����d i%AN�VP~B�ʿf�~����J�l�O�2�P�W��EF�E�g�N��Վ�I��t��Ү\��Z#0{d̖҂���s������&[4��
����� �����9��oR���g���6��?� �?y~�������ǹh}�d��m��V��6�)<��ϴ����"r%��A˦(;�(�OJ�4��=wB�2�ǅ�Ǵ���Tl�>��&W��@8B�@o�	B�����l|(-���h�яZ���1R΄_��N��I�M�O3�m�f�ǈ�G�F�(�|}��ޢSTA$o%�V�8I���V���?k�/� 	��{��Uc��L�E'�4J^�4|��Ksi��h/��+�>XW�|ʲ	���]a#km��ߙ��H���a�d�Rnv1��DR[��>?�O|s��Q�|��6D9����|���C��EB�nL��K*p<�	e�B޶���B�M6�̸ΙN��<d�sR
�ȳr�]-���.|:8��&��Wn���~yR򂐔0���4���9�U����� �zl`֌�?�qq��D�'���d�4Z�E�<t4X�[qz���гh�����8E�5gj���Q4?�tiqǆ�����D`��-K�����_|x�H  �MJo�JIw:�< >8Dljn�.A��va\��d�ƌK�s�VE�i�����b~{p���xj�aB�a'/�$���������co�qU��S���O��%�'ؖ8 �*��s�yW4v���Ck=�ȹ�*l2��Z�)����YrvP�KK��i��|�F��!w��ċø�g����
���w��7��#�(�uu-~),��h������ڑz��7��hX������|�����-�������8��f�8 ��(���ڸ�l�H9m>m��awKJ���]E�د͙��9�����ko'J'��ҁ�A��$�십�A$���<n�:�1)C6jz�͸�a2��b/����v���T$
�Փ%����������*��s��SUU���3@�����_� |�R�[WCD�a}���od[ޱg�Z��Q0�g?%举��ݸra�l�d�}-��5����p�nb��%T�<^;�/6�ag_�@ʖ1oX� �)��pե��m�a �=m��*ϓ��P�u�{�vgN���"J\ �ʜ�{�"7$r�A��^}#g8��#�x�N����n�����Z7���2Gh;�j%F~��/��
��̯�Ǒ�8"���(d6؅x���ؐ�����ht3�A�O� �-w������"��l3�����( �o/.���Q�����ȭ������=�tHɶi��˾qmzg��U�Zg�]�'��o���������u��{��p�2R�X�숐��������N刱����t���< ��h����TI��ڟ�F�<�z�LU��P�!R��'�8�.
��r�v�u e:f��]9��!*�h��ҚZ�������:n������o*�YǺvOjN�Gv:)� �P�x�n~N,�]M�z�K����
�:��7���cS����ˮ��j!���E�h4�G,u���@֓�����ĉ%��'A���8����|ؿ橩�AN5�N�%�窢p�I%�mNS�U"~g�̢��w��=d7��#��u�A���]ݧ3�|��õBt�I��zxj�.@������=#0;�*�,��i��.L��B:�|ht�A5
v�6�|)+�ᅀ����M�q_�X�c�(�1ݹ������eV� �eq���� �@f-�{(s��yq��53�V�h~�grn;�������ng��(�jȎ_f��+�Mx��xN	�Ky��KC������'h�I����4n��+Hqd����3�.n�\yq�菪�]��&�v>~�`�[{�Pv��<�`<�����B�w��4��a��\���Xm
�b쎋	I�G����w�|���+Χ\�zC�Ѧ��d���o/IE��\C� ����5�����s���l����3D�a���~}��{�ފ��O�$�W���g��Q�-�,�i��1@�zf8�Z�DN���Ԏ�/ڢ��"V�!�2���TX�e�TF�/�M�gr���	���o1� 3�A���I��-�����Us��3�PO\��U3)Cb�9|F���y��^bT"��\���w>��� J�!���X�����vT��K`���Fz�]�D� v�y��X��R�7���`���P8��Mh��C����R;\���tE��1��Eۢ}??�S�1���������FK2N9S5�����BiN��3i:T ����iGsц�]��z�����M7���ƚ�!U��U�l֫��l��:��n6�~�%4���v��5W�)T?�%J!�q�m���y/0����?����[d����IҲ�wI�.�e
s������L����I?؂2�+U&R� 1�3�C�Vp3l'��	�OQoÀ3P��X!8����WVm*33ٱ�AM�^5`�J�;��D~���|���U���!�2�R�r1X\,�N�8ʒ��w����nn�QS�o����x�� ��2F�8h;��!�K>����%�bK��r�m7~�G��>�Ѹ��ٱe|�&��K���\��1��.?<v�vE]�b�h��	�(n���^ߙP�&��4�E�D�<�y�x�2�Ώ(��=Ԟ{���3�A�Ɇp�I���5��-��r��ׂ��ލcoW�����'�|Fۻ���S�ΣQ<R/��re���ߎ���V�#���4��f�'����ߕx�0I�^b2�ҫ�vd��Pй�� aX�3�T&�Q��֬������:C׆����[��kO������'r���Z�$k�]B��6�:�"�~��vL�=��z]�A� YWU���[�&
"ɜ<{X[\�m���c���S!cW��C?��2F�.^/|-{#)�J��>YI� ��&��m��1h�=���!��QI6=��2��7��Gf��yn�3R���|���J����8'��5�@���Q(<ŦmItt�-�hH�
�l�/a�֖�I�Q�?��॓��S�|0i�bE-%V��1B��=֝���͈$�@�>g���j�}nC�ctΤ[�dbx��DR}��N�M?YJ���o
ݎt���{�ñ�R(�M��/P�Vk���g�=����I��Dk��7$�A��������D�au8h�vǇk5�v��D�`fK��cJՌQ��B�G<2m�N�H�(���r)��<	��[���S���������1Ķ}\�����	���E��S���u|�O��VD���^���"0Zc�ĝ��<j;q���Z�Ag�wS$`�c[�ě�v����<JcNL�z58���F�5C��jX��:���:}:�)d`�.5Vb�0U�|�Vc�� �X.m�ArL�:{_J	A�;@�la����s����[Y'U��79є�E���M�#�y�G�j>\4Y�W�~K���Ϧ�f}�A�O	�s���k�'Z��]���f���������e���Y*�7]vh�!2Ϟ��@��Z޷@Ɂ�e�n�h.�Qs)B��^ʴ��f��Ր)pp����$�\����Ta�)5�d�v��fY����*d ��$�	U�g��i����M�~��1���94�9�uD��g�桤��(�� �K �Q)���3r�\��%@WR��)�����3"JW�q�~5=����� laD�m����Jx&Z�Y�=O�� ~#R�'Q�=�,��SE{����/vrG��Μ��(r�����O�.� �Z����zAz�Z����ٹ����d��G�Ih�Y����o 	�� �M���SX����r����I*)#P9���Z	)��"%U��r�)Z;�Qrd��	�d�ԽT��e�xu�]��V���I�(0^�i�1��B1 F.���Rez0KΩ�Wt���FIF&]�Ŵ��s�+��5ϔᙱ����|��'o[�v��*Ix��+l�ɲ0O�@�9sIY`�5�l�� �y}7����u������c��D���שA%�{���J��%�|Jʇ�Uڒo-T�8�Z�1�~������i~;�2u�W ��S�a�`��=�5q���Đ�-E:�.`$��"�و�`��⏳Xub{ wH�s���|p8БH����aNL��a[n3�^�t/m����<�9�r#����
�YVO�t4=u+�����kv��`yC~�#RF%�����8���K�4*+�w���m|��(�]�Dݤ��`�l�Fg�,��Vn�G�̛��ea\��xh�V:p=�sJ�Uk~��K�������c����#XN����O��N�wWo���9:����K�M�zj�N�~�i����R��0��O�m���pR��'ɭ�&��ފ:��n��\|�L\�.�L9r�Ӵ�g��
+�.�19^H�f�3z�z� �Z�<�c�-��U��4M�� �w�����v��dk�L�ƣ���b�f��_]*� ��8VC���4Wk��t\���c ���N��Y.!`�a��f5�R8p�ea�?mS �Q;�	�u�
艨����zh�`:�����߆ y��{�?�3��<0�V��E#��(��a	.�Q9j�zh�<�.��EU̡�턖~U�}?���JeӶ���I"���֢Ř�9g�s�2�o���^�/��^U��|1F����CA{���IE��8�X��K���1oʶq�Խ�#o+fe*[���TF�w��4�$��L-n(L%�-�^�	;��to�Y\��v{�}�Ƹ��B�-���������$�P�V�@U��1����f��$8����M�0���.H-C`t�v::�̴��տ���`E�V���gO&]�]H�>��=ְ��HPu�wN���I�I�9��Նj�|�P|pC�+�I+Ew�m-�����kx�Vi�@���n*E���h�u�}�)�ޤ�οr.F���zd	`k�va�7:3�>�=Vh��G/���m��T�2�/��0�g��y��/[HI�j�����MvU&\����d�X}.���E6p�����/�iF���SQ
@99�5������ҐCC�ZbZ(a:�^s��Sj��}p(ؘ�m�w��S~B鉋u� �:�}L=��vv�<��VK��L��������t�%�� X���gg�K9g�CB���3O?`��a�Q�!5��o�Y�7jXk�p��}J����N��Vu%Q�����/�M��*��{B�$�����G��M� /5���l:@�����f�,;v?w���BZ�x����-�A���J_[��g��ݵ$��%cxm'�M�W�&j�֠%�t�ZH����(����4�D�>� �d����`EEeK@s��t�#��z&�?_/cr�<1�$/�+���P�E>��0|� x7a�e�P�٭ec�e}Y�a`kX��4��%�֟I ��+:�W�bw��]���D�k^to�V���hP��.#�9IY�O�ʛ�H.�`�n��rF�f�i�L�I�%{v��?�������N�=���,���B�̑q���K�:�|j���g�mT�b��5�ù��I7�L+n ���<I,�u]���~H�`���q<���X�u�)g�.>yv��W�M����ePU3g�-�3�Qe[����t��]��� _Ã�=e��{^�,�c��T���R�����0�.6=�2�~`�?5�sF2ç�vb�ͬAZ3��I!UX0$��kҌ/i�O��{�L�fR)����z1;b�v�!*L,�v�'\�A~�!m(m���.�<�����@�ъ0��?���
V�5PTՅd2��``j��،��<����J���h��G/�g��x��2u�g���jFQs�8{���;�_�h�g<�셁�N�����L���`]�CuT��9�B�ޱ@�=����O?�`�i����Cg�2Y�"=��+rZ�hDPi7x����I,R���Z3�VG.���H�!*�'B2ƍ^k)�c�{��AԶ'���l�Z0	��I���Y��WхFe��stL�R�I�b���s��Uf���13�#fS��x� R{�pȡ�dr(t����OxY��L�>��(a�O�Q��Ğ\j�J��*�#��jYZt�7Z�ԼP�+����t ����\�ţ/=Ȯ^OK�di)ͺ �s���Ҧ�M$�Y;`pؗ�ml:�
��& �!�W�xM���ڦt�e��lg�Z�v8Tʈ��'o�A#���
�_&��̱�{j[b��Z�
��+�rO����m�_�s�'~���Ë����k�����޲�<a�"��L� �X�۽�Pl�N���J���_z���'e���K�\�s�ݡ���6�j���w�8���Ҏ�d�����1�⳵�Wc�āq�lv6�	B�	z��0o
V_�96m�m�E��]�j�ΡO���w�@2�4�@m�(/�o�⁣<{��*���T���r�+��2�&�iWI�k~{&�1- x�Ԫ�P1]���1D���m�ʕQ҇��a�z7���}F����p�C�ʏ�Fk��M���G���[��[��v��!r8���@_cV��[^Џ0�ۡ�����ƾi$'b�����pB�?�%,��8��_�� 5݂&z��	���--��r���hn�#NU\�_`Y)I������_�b�F�̺(*��ԣ���6*�U����I�h�Y58N�v�rg��tۇ�����9(Փ�6�;��hi(m�p�V��dOc�2+��:�3�^�%���5L��ա�R�-Da�M�];HX���T�<�����j�5�2��(�~8��U�>6�Z�����4�|��l�x�_Ơ�!%�^PQj+V���?������ʚ��K��
�z@���%;??Vh���f{ح*i�[�o;)U.�&A=6��Lf�/.���Zi���E#��-�u�8����W1�Ծ��
�Ws¸zr���ݰ����3����aH_�|�Au��_\����d���N	��VHR�w#��UǠ�H�){2v���;99ݔ�d�hi&��_�׶,e��%�8��)`m3�X���S���vQ(��۳6��-�CL8="�;�*� ��Md��s�gx����/��q ���s��x��(�c_4����^���}Je%��2�gԟ�1=���axZ#��C�=����������gn���x�($���B���feHKp,�ph�G��Oݧ�C���r��\=�hNsCփ���� �w�Ձ��
�[�o&G~��-�h4�gҼ�E>(�� �+�m����%�(��}d��H�����D�]0���c����)���o��|6)"V�9�CEu�!k6z*�/@?��M��K`aGU;`S�$6�b�9m��V��3��~Y�A�Ȫ�N���?�1�4Tu=���7h��?9���M�Pl��x��Z��'[�Y+^�c����L(�o���Z��0p��҈өsTOb
j49_�|�#�a����Ĳ�E�$�:[ԕ�UG��K2v`�9�j̐P��E��p�&wJO
�dd<-��!*t�����-�����QyJ!�
)����=[F���Y�F����km��^�op�b��� ��<��hq����k4*,՚B�d%(t�O�E�I��ʯh�h#�7,�s� j7�U��u&It�'u'��=�ح4%��E���m��(��,o���y��ˋ�|nnp�ci[���������c�z���ܜAT��E�X[#�I� �z"^L��׏0Q?�^��aR��'pD�y��Dc%����k�!�w�Wޙ�nt�i�B�t���u�z��PK��`p�خ5|ލ�8Å��^�:Ys��aq���Zi�v.��;�&�0�4d.�����o`�q�]Y��Z`����<�o��%:��f��^(t�ዪ��;xOǯp���VcWO��7
	������	j|hwQ��P�U��燊�j��в|�N�6�3��w��5��&�����_�Gi=N�Z3�E�qF�a��|��_���끚lh���~|��n��"P�}lG�&
�	c ��_�3�ASp����`��D!�?��V��ࣱ�X��}����Ը���-;��l��b�^0��y���oМgiX��Jg3P��ςB��R)����h��IR�JP�@ﴽ���.Vh8r������Y�u\�.�]FLaڂ��b3��&APzȽӴᐵ�F��������B�~�o�`��+��������� �*$��G���U�0���bK�j)�d�9ו�93�B@�	=+f�H��/��^�.3ie�?XJX�+H�wi��d�d_ޔ>5���;|J�+�evP�yRK��a���b�P�?�;�9�J���*�CsC��GL��M�׾�n��TJ�&�e6�����.Rh��ɌptLx�S����J�+.ppU֌)�7�I	� 'C���b���f�!J]{%�{O�P���
ϋU�K���%a�S�������B��5���kֹ��̈�Y��z��l1��^?�P�b�=}�o�T�בg���l��m�ؾ�>Z�Dw�&AX
:6+�f m�P�x�|M��v�,����ś�/t�u����$�k|�sB^J���z�OLiW��m��u���뒒�}���N����&�X8-/$�F���c���v:{o�h!��3.d���t�g�\$�L0;�������7��T�W�/`�@�1�����(����$������p��`(�'��
|��!�',�;<H�6��η&�LฟZa��+X�XȢPxH��P`2T���*Y��8��n��Gu;S�E������{S,����9��[�A��`߈��I�|�첼%��?f3^#��ꆂ�>&F��-������C�}9(��(������v(*���(�;3.�`�S�L��b騨�^��I���q��0-�����*��ð��(Ԟ!�@#U�X������TY�U3t��`�� �ـ�;�c�K�a�Ȱ�fP���h���RD�q:��CDC��f�M�D�=�J������A<P�Z�w�AN� ��J�MVq��+͌	�+A����ebW
a��l�OB���>ɣ�}����}0ũ�h5�?�H�a!)����@������9�����oLY��H;��$���a����VF!燫��?�o� 'G�����|��G���U���d�\��P����B�~pT"^���}��$���X���ah�6�3@7ɖ��*���x�A�F�4���&]#���*��Q,�^��2yW��Y �}��S3\���rbk�j�Ă#Q����
���*S��<�eϭ?
��Հ���u�Y�]��-z��G��}Qr�hQ�=�uo��τ������**8���t=uy�3./�щ�y<5
6~j;'��s?A���TRU4C��Xj�/� F��tԫ���s=h�%��|��T��w9����G���RrK��jh	j�F�_�������ޞN�U!��s��\���M�x(���r:.��7�h~�(�{RAR��d��v�Z(���Ϝ���j�bjp�ތu�7�0끯d=~x�EM)��Xs��JkIJ��+S�ލ���u��;���l�-A�d�&�O٩̊
�F`u3mo?V�i�>����!U�|a�͓�[i�uS)�vA���kç����q�\X�7�_�n��5O�ƾ����yp�ڵVL#(c���ds����C��O .��zB6(LdG
����Tȗ�@5+��+�.�0�Y�vϑ���
3���b�yW]&W�O׀�ó�A��eCjs���n_�pЀZ��6cnG#�.Z�_�8U�+\��+Ɯ̚6�}7kS��M�󕻎��BcȲ�Շ�:�k11�se��C������1���,0WM�G\ ��ｳ8G���YOw��.�L�>?YU I-N�H&҅���<u��W�	���Ͽ,���W0�4艦���塒Û5H7�d�C��6-	=��\Wl`
�W��`�]p=�j�TֱRm�X��3�m�s_G���@w�\��l\ad�NU;���Ä�)��cj7��s��@(iT��Zl��	$�*H�޼zݥ'9=��3��y*(s���~��%�-���l"�w1(�ˌ���3))ua&�'ǯ�~w`S���	��آ ��$.�;}0{O�C�U(�Xc:H��W�.C�3ߩ���/��x�;�gJK,]�)`b2k*�G�ӜLs���@�A��]L�ƪ�֞Jf�֚�䭎CriP���@����
I���Y�7�7"�S�(Nht�
g�e����-%���>z�)%��}�_��������	rJ mny �U��e����Q��#�&���0��"Z^d^6v.M )����_Ba�H\��_�i�����W�-���:.�ytEY��<
���5�i^4�h][�YYF��JIp���1.��(�.��J����ħ���P+���	BK)`���=�B?�3�i+���%F��5F}�w����F�KYgUZ�`'ɹ�ӆ8�ɬx�S}�;f[1�Dw{�s�e�f����T�vB���~&ΩB��(�C85
�}Ld�m�cuQ��)����._:����z��6%�]�k��,����\�j����7v)��c:N�����*��y̻4<8 Ϋ�&p45���X���1�ǚ����Iy���t"����^A�����n��ȋg%:�K��x��%�OY�\�<8_3�%sI��]~����E��#M�;��n���5�Id��i���pS�'P�J�`���vmmP�Ҿ�B	�p)ZNN ��Nc<�[4�A2-a���:�]؉�2����˦K!s#�������f�V����D���)���؛f� ���'�'u�%�2(�Z��t���-�< !���"ڢ��R�=.h�M^�^^����>᜖9�]DUl=`J}tr�*��\?���y!h�����Q����1s�L��(L�ҟeP�7�ĝ���~j��1�������[V� �Z!��c$�q���%�������x�ncN�A8���#Ŧ�J��[�_nݛyPk�S�^���X@�ǨE�P��^���(s��V.n��I؂G��B�����:�=��St�`�]����/ө�bZzX�9�ac�FQ,�C�Dxh<D��,��-��x�<��}���~��'�UO�H·��_��A>t��eμ#��)x)lO�wsߍ�N��4��R���b\�~��m��i�sr@AжPt2Ì��gT��o�۶�a�I$%�A��=5�Kwꊂ6pE`��Vo�.0��L�t� @���C�;�&\���*�l�̃�w4M��VP��d'?�)4����Oo�u�J�lp��P���4��� �L�R� x���rpI<������I_������Ͷn%�`
e��,�&�;?���\e�m�F~��6���]��f�3�~S�	Ҷ�7�Ǜ5������~nST�:����G��0��r��X�oS�c��`�n�a|�L~�՘��L�:p���,�������l���K�a��Rg]�e��bu�r𞂇tiE��-�`���K�I���*u�T�#!�����=�g%`�Q4ɦc_�݊Li�T�	X�E`�g���_�ވ�������%#sz0��~38�0ۍ��Y^z㏷p�_�< ���	1O�X=m��m���6ĵOM���lv����w�@��,Ԯ���;p�¨�#�{s�s���[F�,�:��-�f^P�BFaX�{cVv�����;���/���^G����?��$��u�`�+�zrb�э,Oke�^�D��/�#k+Q���'^SF�,W?��_~mXV���	ؗ�$糬�~	�o��HISl�ۘ�m}R�V�ʞ����gh�U SF,�Q}X$�5/K�⛵�7�zl�.*�p�۵%в����h~��a�f6�ಐT&?��r�|R�lg@��wj��`��4>{������E�X�}��0 ]� �y'_k��5.*	���9{�N�i����rz`e^�s��ӿ��YO��7��b� �~��u��Z8#|uY*�0u�G��s�f�[nÈO0|������z ��Ia�{F>�R��O�nh9�4VwU.�G����]d7pi�|�bhRZ���7즠[������)����ưÀ�)$��_��To�mؾdr��l,k,�~\�`������5�5A��.~ʚ9�����RT.���7d1:�db�0y��ũ"(c�U�M��㯺<��8��Qͼ�#l��/��	J�喢�:]�n�{*��B ��l�����Ϧ�q�v�e)�G��րb='�hZl3\�1S��vs�J���c�Iq� #�X���c+���HwU4B��eG���Z>V̴D�c+ڲ+�rk��ቊ[Y��5$�l[����vt�k���"he�&C#w�DqE^l����'.)�3@8m�[e��ZfH,�3x���u����]��?<G��V�\�{y��螠��ᇂ�bߥ�V�p9B��c.$b/��W�.�	^�}��_b���_Qu�S4�C�R2ײ�be�g�âg:�p�IϚ?�\)����V�Wlяr��yá��'=�{�e{�>�'�Mb�T^���36�Ze��)�f1�XԱ��j�̣H��sy*s3y'v�Td��k��%��?Ǽ��7��	��8�έa��T�_ҧ���3��| s�AI����k�C�V��VZ���t`K��q8�c�k�����W�(/P7Y�ɓy�E�'�L�v�CtD	;���{����� GX`C��w���~{��ΒH/���ܣ5D�%oѲ#�ml/�"gv�hQF��/i=k��ҫS����:f���^
{jNL�$a���"纄I���.1�s���[���������B�nb�2�!�nUg=6�F�n�%��V���s�`Â����{��
}�߰f<�<EY�����P������U~Q�����.\��j�he͖iP�-pk[��)JM�ހ9A��!a�o?����"l��cu~<Ɍex4��#��AѼ#�nׄ��b���X�u��΢k�ߘ_w�P�]���i��Je*-HHAI�Nb��+]�7<�}�'0���~Ni�בٵ>�#�
�3�m�5����%�)K9��A�@�`x9�B�%Imb��=�T'+h�j;D�q]E(���DF�H5��ͩ�k��z���F�/@��iMs.p��`4�*D^�%tؗ�ͽ_�1$)�.��5��loW^�3�W�Fv��X�`�_!q����3����8�p"�ٲ�F�(w��to/��H���p�} �X0�2?��ȩ�����O�Όf�3��StW�46�y��A�BO��>��Q�K�V�A�)���j?�Ia��/��.��͡Y����"c��2!�@w�/%U�k������?%���4*�	� -;��n�S��2�������_lخ� ��ڞ3�|�H?=!��R0`etIu���?kO3�rX�
ԁj��ǈz���E�rTsq��G��\�M���n��#��^1�Z?�@�S)l���@�r�"?��L%����~���-�)�{�f�zN�b?f�ǬpB�̃��@�m�e%��-��x�������E�v鮰�!r�A{������q��l��V�C�Q���k&����	�Xp}��]�AN�����.�M�b�r�~l��f�x\�5��XN�~�#�a�[�g���?}]ʾ� �HbZ�J4�[+A���³�>��['��c�mpx����� �zØ�TH�|��(?gnv��]Zsu@'m�*(?�Q�����,a:�_��z��#{zy2��_�_>�ڍh*DHϦ�gJM���)�W��g;���r;�ǩXY�I�Q�x�B�cQ��kW�o�)f̞J���"�2�\���je��z8kCl�W���@����|��u�I+JT�p�2��~�Eԑ��k�θ�޿Z\��~́ܡ��;��VⲰ�cc�I���Na,�u�%T���*�zNJ�5!���u|�y��3s|�M���٘�zv�����I���P\5����#��!�$P�(���ZsP���⍕���q�$ݭ�+
� Z�3lJ�  ��� v-��$��tՕ�����9����W�:'�<���ќG��k!@��-������*m��?o��I5�֡��c�r�@x!�~��?���`�V+��ɔ�� �l��7��/���(a	t#z�����͐�譴�u$�S�N+%�l�B���9�h�F_�J//�q�`KV%�;+@K��nl ��$��Ö:lE��f17ik3M��k�.�ͻ��)^_=����1��0�,2R�\E�=�ڈ���V4h�K2�W�$�9�7T��Ѣ����f�K�w<�!j�ܪNm׌#}�gh�n.mp5�@<��2��K����M��A"L��N�gSӈ��$�r�TY���^,���(6v��@7���F-FK®�͒#�HG��V�F�c}�}����t�#z8���w��	�9��5�:;:�_��0�M,�%� ��,�|S�EmyQa�	I�Q��P��©�k@&,�nj�)���%�*��̳3�cs�8;�4Ѳҁ��0UI��0�����e���2|���]YI������[DGY�n��7k'��� �E�wP���/E"W֐]��Vى�]��,ܲ�W�z���i��v��U�� �	۹u0�.=�����v�1?��3�@�ӅG��@�	ˊ�x���>��GVq`��,��*Da^�t�V�����Ԛ,#�I'�dN\����=�&��k's�P�_�C^K����x,\��Ru�.���8�/;��Js�p~!��s<gctkl{�.4g�5j�;�zN*:�Be�����|֦~P��N���G��0B.�������>%'�R�n�c�W@�Fm�G���_D>��������<��,9&&3�U�Gu�1N(�g����ob�oPJ�Rh�]�E�ٶC���:��+4��%�����[Q:
ÚT;�s�p���H��k��_�$�׳��L�\��ꅃ�|G�ݸQ�WVrr͓:���o]�B���jvVAp�hp�����n{�<�Q����?L� ������+���?-Mwe��먻�~�㵕	�)<WS�UN��	x�i��'��5�	����ū��,�( QP���j��|�vN�ǳ5�L��½	��m�t�4P��H֦�ĠI�Ft�4�啄D�5偷&������P�1��	� M�ի�-t����<t�&������A}#B�S��\�����ᘳ3s������V��6�� ���\v��a�|�u���&y�kҹy�t�{�����0��:��Ȼ�þ;��=n�� Xb���������)$��a����ͮ#�i��^� $��R@m���F�����nXg�֞͒�R���Af�
O���t$y��1�ѷ�S�j���]4��:�p��)Yd��f�OL߱F�H��of�����2�j/���@p$�,VxF��)��b*�ZI�� r�o��gm^�O�aY�dA52]y֐m�
vh%>��#��:h�����Qן*�[�u�e0`���PٮY�u����� .�:�/O& �A6-��\fk���9�����?���M�xnqq�D]��*��n��~{��9�xs�
Q�6S�O#KE�������@%.s�
��/�P�����E��:���6����i��z���0��՛�s��7l��r�8��L��n�f��c���'ч�����E��>px_��O�H|'#c�a�w���� Y�j�h�<<���绠���<m�S�-3�k,��Hd^%��\��nc�*�ܲ+R������d����V]-�H	�7>�M��f:�Y�m�d�E�j/`<�ꏦ	�������F�ަ��d�F ��\�}"�=�W�ͫQq��`�/��v��כ�Ӣ���P���+X�c@�`�~aАk�Е;\޳�P������f���Z9=Y����$P�k��6uPr�=}�0yL�-���"ְrN�R	%�A
zs��;c��^
�o�-�C� ւ=�XQ��?̉��$`�ȏ7augh������t��S�J�.�I7�$'C��/Ij%陥���6�dzN�=�+��y{-�BA���R�pq)�	���p�`���B�1�F���}����Q_'t�II/(�ղ��=Kn�j���+���ZIH�,�O�8,rV�&�hғ�ׇ�Z���u
>�3"Dh�$b��Hّ")�='b\�嘿�M:al����;Z���Ʃ�5�BkV�U��<��w)����Ƃ%�0�����s#���
�޲�&���[��Q��>y������yvzQݸ��tbn�iiP!�m��|��~���W/�(���
�n�\�#-U���+�H��-�W��@�\T�oɉ��-L���
���8�'Q�`�?$><���'"�ħM3�	;A|�QRx�|(��D����D�ĻʥР<�92>�t����8ݴѿ����3O���*U�Uq^��|�
`�p}�׏]��g����ٸ
�v���{D��RT��1���*t�D;�kM^˜�A�"�+�%�_�Ѱ�:�0P�h+�:�A�gٜ�Ï���N3B�m���ؐ�%����n�����I��=�v�c>L6�밅\�Mh�
0[��'�������U�K��YO="�0V�0���ϱZQ����AVI���q�.��9��}�7����7��/�R�N̛2s$�F�Ĳ��� �1�b��$~��?��
�g���0w���2L��5j����Q�uL�Δ�^7W�7ב�~3I�	Uq�1TL�gf��s�p�JpG��6�a���0J�F)&�s9�э���=����&�	��z1�Oi�z�]��{�o�;�{k	��W��tG�IH�2�ÿ��).��������u�����\�6�8�W&M��$�GA5Ę&��}�(q�9S��1�Q�	����T��[H�d��~��JB�ue��?��)�Y��t$��*���>�g�TrL�#*�5L����<�0N�'�B%���"F� mM�`܆�:a4f]�I+�KCH�|:U9������W�_�&v�|ݴV�1�@s&`�ݸ��kxO�S'�Č�<��-�Rǰ��*�5M�*�9hۮ>��L�|}"鿚d�נ���
b��}q�EL9� w4���|������r�[��@�M��ޔN>lQmC�'6��8���J�¥(��:����~�m9v�ۍ&��`�md��]%�_?J����ƒy�W��ܘaWD�v�S'Kck���a���ok�l@A�.O�� ��=m��;�^����eloQ�ާɦݟ��6�\�)���ק76�)��K�l�j�nG�`i��ŻLƟwUa��i�0D+�U�X�o�1��$=���i�p 8�P� ��_!m~v��R�4M v�8/��%��`�ٍ���<+�o�ߎ�8�����(�I�D8Y*�:}@,�h�����5�t{鈽�}��� kH��<�\r�?��K]"��r�w�r�dx6�ӯA�r����Y��?�;�'���t�������ɛ�(1��Y8@����6�C�e/���92&��󙢞m�����my��p�����Y�pZ�%iA2N�z:�A��Fʞ3KnIPy�c|jp�J@X�-���4"R�J8K���X�Rq�����"nI}��8���#���s�7E�Y�!��0Q�&t�no��-ע�	'�ZBa��͔`��}]N��S3����8��<8d뗧#Sy��� B�m�H�����DY%+�d�z��C ����^ڄ_��3�ڼ�Vd"��Y 
�p�6;5�)*'s�炙�nh��1z�#v ��n.��B+�w��x��P���ڶ�"8 �5�J�ޛ�����A�2ʯ�E��j:����Za��{�j�UN� �2��j���\�ň�����(Ȉ��]H��I��&ok�
m�I�]�'�!�
�_�~�lR�>"뱦���$f����f3�fPf�[ȹ��z�#������/��~~_��}�E;]�O�/�Y���nl�~��#P�-�M���&)y�����t
�3����������7>r��2�o�.��M(� H�8TY=� XY�d�~��Z���<p���[�tƈ�	V>ϰ�����}�s��3����̭���f�0ұ��#��95f��_�ݹ�w�UFH�鹔�H�P��';*E&��9�k�o���鑥���b-��m6,T�D	�)��B[C��&\��P��c��a�=ܾ���n�B�(P ����2Y�s}�����0�<�#���2� V*�/�>��*�A�������9E�.���� �w*�g&l������Qc\)��5r�����V�6�4*mE3�%���Lߌ���W���J�M5U��=}Í0tb)@�zkh���"�Z���f�kӭM�
ʱWl� f��fŠ ΩYh֭5� ��b��_�n��@�$������6���N<Q������nω���;��t������d�A��M��*��EN��2��Ź�����,�R�ڕ���a�Mw3"u��F�V�N����-l
���'�w�!V�exy�U�>�	*�SM�3�Ӑ�԰�ܐ���%�)������d��>����>��_}?lv�z��a'
�}dv�}n짓%�$B��~:m�9[z�g�K{(Yv�����+K.�l�ܓ 
��������3�t�,���Ѽ�እ]�tݿ�+"�5���O�P�n@=��/�e������G��d淒懶t9ϧC����ԭ�'s9�n;�g�d9��@4�:R�N��Jhb)}নՌ�zeS�'�<���,۠A��J�6(7��F	*�����bH�N0K�ʵ�׻$�G�V��Y5��i_�&:ia��䕇0.��&UR�NC$����j�!���9",�/Pdu�pl�]��l���;|��}T�K<��)�c� �Q��E!�kO�7�%>��~��f�1��d�-�C%�^��3 {q�A�&�-*�|���Ń4��kP�}��Yc�~"8B���yf�j��?r}�܅���?��Oy6�e�ύt3>�h�lB��ɔq�CHR��ȳ��X=�f]��[Ո�\`޵"#�d8NW�q#f"��t7Z�|�0�TN�P��֯k8$�L�V ^6;�S��47���S�k�6PhpX����]��R>&����B�'�����T��>��D��d-O���GC~�jhE�s����`�H����?4a� 笼���|Vw������ą)f>�T��M��CBu1�6�w�B��-���0A����*��$���+G�O��n��3���XH����0h�zϴ�	���I�%y�_��6�!����"�_�p� �l�r��m3h�O�X�5W��b�]N&��֦���}.F�q�`�o;���=):آ�?+޶�U�T�r;���Ϥ�@����3;�.]-�v��o����^�Ƀq�ٮ~K�.�
�3���/�̈́�43p��2ն؆��3d5���:������B���@�^?{څ�Ԥ�I��ƒɧ},���^����>�����q}<9��t����*h�Y�A��Oפ�����5��n��A�ܖ5aYi<�L���|QfZ�G��тh۔,N�e<-���cѬ� "��>9&�|�>{%˺�_ҫ":v����t �ߦ���/���]��%��:�����Z��+ڐ�,u�EZ��?�����]��I}��uQљ/��#������l��4Tʳ�Bv�Hi�V �Cv"��(S-{��i?���Fu�#����c���/�鯏����*J�J\�V GOU�K$����N<�ю�[H矇F�S�L|�g�O�l�[ӭ�_.X��E)�y4VbO���q��}-X�<��	��*��Ӥ0W���ژH�˹��+(�E�$bh��P�z�~�1K��C'��^�T�B�wS�C�\S6���Z8�l�gd*)��n�����t̨�η<J��C�����(���`��а����[���;�1��᳸�{k�<Kq&*4���ˡp�&�5CU�Ƶ�pEށ"�Z:ݚ��h{�Ù磤y�1��2FBi�I��?��e|KH����LC��/揜]d$�k�m���F0�����R�=�>b�hF/��l��������n�� �go�E�����&�I�ӃN�v��0��L���1M�D)\ä킬��q��:�ő�'+�)�e4�d{�����N/u��o��+�̉��݂���S;C�& ��_�o��=˟�6,O�"���2șT�ŧϚC�'�
h����T��0�;�QX೦~�������K|��ƴ�Vx3I��C�4uOR��Q�;���1!�;7ȩbW���-LTC���{��M$���a��1HY�u���W���X�q��|��[��IYc��)�e(�,-�L�Y5�*s�V"��p:M��T�64^�Ow��OZk�\G��n���C��:��I�L��X���L��:o���hi�-�V����-���!�� $�4����1~W����>Y�I�^kD��:������Ե\�y��Z�ihH~�f�I�ϫLz�)u�ު���i���&7&e�w�� ��u�����<?����lfXmV����Gp+��6�������br!lA����U.�(x�M� 3)��m� ��q�~������������ț��	⹨X����K�1?iި@}���lb��Z��*(̤G�%ܸ)5������ܠO[7:_2�c��Ж�rIje"��Wn��c[����s͔K����~k�z��R[��\�=�� ��t�����2��U$/�x2%s�[YOI3��p���GV�1�W�R6|뛇4�|*I����߁��~���`�y=u\o��C���S3�/��Ǻm����9 �J�k��V��W��8���1LI�a���6���-S=4DxFß�� �"/%�t�ҙ�����ŵኁjS�ID#��1n�!����2�^.�����Y̩"0�U�:��v���lg[e��J�}�׉�>��
%tU�Y��M�ɢG~)S��A#w���Ş�M��9H 1���aB��E���t��K	�S�����N�>�Ϧ���K��L����[&�ʊȨ�-=���#V�T��z\g�@�8]����ף"Ҏ ��N(���փ��h�cP��Zn����nA̽(B�΢V�v��-}��%�JV��sM�̾�a_��hS=ier��'c��%��,a�<ߴnf���sg��[�W��3x�oT9�n�e����+����`ԩ�9����;�V�:�	#L�F�!C�ɒ�b��3v4&鏣oD&�W�%N��B�L�	�e^�Ζ��C1 X˹��V@�j)����O�X�{��4���S�5�Y�ݦg���a_��jz��#��ﹱD,	�COژ�I6�DE�MV�	�@�hDJ(Г�m�u9��O�������SN���n��/2��ZzZ���%6�W�
�1nX7tj�?���$���$���)�ʴr8�A˗
Ǽ�p�.���6���ݜd�'{J׹/F���Ɣ�&�E�bUq�`��KJ����|کաa3�b,3���DE��Fo*�W�C�	0��[
e�	Z��ڞ`���fN¸2�SeSFQ�I�ݰD@_�)U�`�#��~���$"��/R[����Q�'�f�d�ͯX�[�)�����(A8-�-
�6*�a�����h��~�ʋ˙=$��%�j�7{��CZ�������{�@4I����є��jiR�Z�?����6,:P�JQi����8��N`���Ƥ��ӥ��>ɝv�|985�\D-/t����TX�l��ϴ��j!Z���_L�"�x�'
g ��X�"�t��r�c�R����	߀MSk����J|�* �)�}�v�G�­�k����&��¯��YP�A�[zS�u�$5?,Sq��z_,�9��������J&>������hƗw(���vD���s��	{���?����X�'�
�t/g����'�Ld���ZFbI��>���t�5X��s��6�Ԭ%SBi�7�鏙��4y\���`���6F(ji��+�G���x��x-#�n2S�|�F2��#>���/�.��Qd��Юy"_�Й0�=B2RN� ���ۻ���A�3��^Wf{�Ul	��xM�M��۟���ed�=�i�b��P²Z��멱Tg	r� g�S�Y7:�N��Uj��;a����8`��#\�����\ CY|Џ�v� �q�MRRt0�9�G�S�|w=�A�������9�i��P%*�C(��u1B�G"!���,VU��mΰ�ߘ~�n�&eP��~n�����L$�h"�OJ��5��j�i��Cw�/1"�//�?V-��<�PZJN@�� ��G�!��oqC�����Gw0�r�ja��L<��N���ӏ��#��DJ�Sd��W���)Ӫ��hըLO���9�+���S�š�S>��`Zl���T� ꡃ�q�<tR?=�>�7���$(RY#J�e@����W�a��UB��W �ڈ�4vGǢ�L�7�qJ[Qş�	7�=�}.3��'�{~�M�������%��r(�i��K����'����)���2X�X�<W�'��;�F�H31m;�ܹ��\�v��>⾦B�"�xP�'���^����CViN�ÿ p��v��L\m��ҋT��ͩ߄dQ=����m�����p�}?לc�>�9�X�R����aWEE�� 2(n:��1�Ԡ��|?.vX�"�0�ܑ4���f_���+���1���CT@���`s5bH.�W��rK�`ǨjA�_�[��2������p�J`ba����dH|�o_���~����w=�#����K����8�i��7�6U�D��m�D�'l����}n�U���Q��H���CI��c�f$�p%;fm��n���iSv q0w� �[���CaU�%`<�t�w����`<۠��l�$�-�!� �k�ѝe��?ַ߯b��<��7X�-';�Ճ�I)Ӛ�Ar�$ N��@�b�@p,���~8Z�T6��@;'{k�2��l��e���"�v#CV|i�ʆ#�J��q���k�x��=�=�KZmӸea^s�����Cd(=P���Gs���8�U���LR7T�0��4��'v��OMnk�}��U���e�B�@@6|,�ը��d��b����fHm�B��j����
�ފ��u�?���y�<M��׻
��fx�J�ZV@ˇP���lq}�����j�����4�p
�?���dɑ<w��@d������J���zx0���2j4F ��g�N����qfֹe��'��6b�����WH����<�ԩ���&C��?5�L#��_?�L,� �aC��� ��Ʃ��#E�:�d� �C��z!-ߖ#�k~CPJ����z��1*��g�]~�O�nI`�_�������@\+��N0������N5/u����Z�ٺX�;-����'�+^�&�r��;����S[����Nʞ�j��rȥ��U��B/;�7����d���2=�������H!�5�[��!�!Uݸ�)�^Gи���}m��Nycݦ��CQ����3Af{~�]�2!v<���O��>#|!y���b6[�Y���u98�=�3d�!"�'#`ZJ��l'l!��n��n�TD�Z�9��-������<cx}B���ư7�E�/:�-t���w�;Y���+�燵=n�W�!/��w�����w�<.!��} �UO��̿q)ް��t|��7��Ba`ZkQW��d�É�G魬�)4����Ss�uy��K!�)k\`��}+C`E����5q�?a*���`3�_m(�\�a��}Y��u �,��~��P�_y9�?p�/�_�y�X������m��N���cm;C~�r$��$��C�&�Oi�9L���3��Q���r-x�
Z��2�p�Yah�K+�"E6Q�GR��c�����l������F��O��]z�vsx��v��B��a�0�������ߘf�t`�?~Q���U��d4�U�.�s��NG�VZn?����SRP�Ǜx�«D<�J��fzOTzv��,,��;u��u�ez=��c���ń��/��S�L{�A���kx��G;+���bE��IiS�l����(	/���Y�<{�3��F�.6�m������g����$�K,�����1^��Wե�U x�~քB"X��9���ݲ�1Q�����L����f�+prsyM����Z�/�s+��I#��J���r���6�8%K��9�n�;��-��1s�e�U����mge�y�fT�R�!D֪�.6�_	>��G��*~Q;w}5J�]�=����K�4��Ǒ��Q��笆�`ϐN���/��1��p;)ϟ���Z�3$����Q��R"�N���pM��8�@��I,��W��W��Nl5�W�)���&I��,�lAv��&q���ށ,�u�t(�1I타|>9��r}�ˬ���a��(�r���5�Ë�˱���Pxګ;8�<�j��Hv������]�[d���GΜ��]10��4�;ӿeC��/��Uu���vR.Q����c�#�Րҳ�ɀ�m������^�>����9��h0�hSua+�) �	6¿� �Z����揄Rd8e%�+��*��s�陟��^|,�-D`ZIQD�9j���fx�rht��k�fqY�˥)Y{<%�j7D�w8w��SU2D#4�7��$���.�f��b�/0���Ot�!��D9!��y�9��7��BF��fi��̯E�:�K!����"Ս�o9A�Q��p���)6�;�1,ⴈ*���y�vʖխ��]l�d]N�40(���8���0%q�u��t�7��j�J/x�A���3'x�����EQ��no�,�P�
r,��2��O:X�z�1#� ,�$i5o�ʜ��9 �E C[�n[��'�rZj��O�5H�7Q�Z)���:�]|A1�ܲ�6~�V߬-��U���xkp�[h�h�Q��Wc<������V���p�+O�Sn��!x�d��C�`%��υ�:7�گ	�Sv��ގ�C1��9<���O��aH6�Mu�P�&'�'D~յ��J�Y���-AEl�E$��v�l�,BFFQ%5@,������.� �pǟ�]X��u�7����|�aP�%����E����
4���(�N���	�T���l�y����{�˗���Ek���A%jb4r���⑹��7`����	�#��E�7J��ؖV�'��ᷡ�RŹ����/(S�����
���>G]�^^�c��p�S;L/��G~<�������A����"���{Ș��$��^v��0�n��aU���{C�����S�;M�̿r�j�D�]O[B����ӝz4��X4��h��Wc#�����8�Z~��=��W>{��?��P�"aߪ
�]���g7,I�I:�sz�3�P_�*,l��^${&��V�9�TҜ�u\@�?7^��e�&T�t�vS5ط�����~��=��
lP����޵�'$�nB�~��,���&T3`^�q�=�l���~Pf~eЀ6e�A;�Z��_t7�����Vv'��0��P�^�����Ѣ�6K�/�E
����	 w��$���hu'�t�Vc���8)@�54s��5J�
��Y3�\�GO��+W�uҰ�12g��ҡ�~#�gڛ�hp��3"���fϺ��k�~�5NZ��2�	�#Ԟ�X<�{�D��-�b8χ8�������H�O�(�f�T ���~B���R6���5_�`,ˑ.����eY��.V�����h���)=�h�i����&��"(�D����}�?�\�_P|f�K8D�i["~aqsZe�����Z��w��*��G��=Ŷ��/QMH�;}���ؤ����z�LM+	�+��G(�{7����A�Y�+y�r�Q�����`+[,K(��V-�}6z�# .��Џ��E�T�����>̨V�>ɒ�N|l�#�Yg���20M�>$�%W����7%BUĺ�&�g}	W�&!�<�[���>$�U�w~�P5ɔ��_i"'w�N~����<oaUZ�@R5��9�qU�I��O�@���afk�O���ԩ!�AO��n��ʺ3��'���@�������m�س��y�v���qx�D�ǡyS��=���W!���̼�<���1��#*��s��㟴�S'$W m����Vg�B.),,��(Y�Z�942�
�6�������`@�A	ԁgW�w��')�nf�P�:�Ĥf�G��tbN�la�����3���p(\,C�<p�Qۣ�$�̘��I��I��v"��y�Jc_�_��϶�r�2Ԅ��3�y*���'u,C",w�(ϣ�!��R���"���0���4ARV��W,y���SJ����b>�;��ܪ�c-�|����$W���3Fn�����K[aѸ��^&y3_|\X����8j������?p����Y�5�˻��uC�YF�hb�5���x���.#�(�a1L�	}��9?�dIw������52�c��.=2��~�#gF�,�tF	��@!���R,��+��٢�p֣&�B�%��/$��l��BS�n�_5��i�y�;X�ï,���En����Ls�yk���c���C����#���^��+�B�"v�D�E���2?Cv;�$y�J/��C]��R�v��<|�H�U7V"��skP:�7�2�����H��
��-��:+u���N3���ehgm�D��|V�9�_��z�G���<Qp���/m�i����t�z�u9�s�����?)jN#���2}��ay#ҫ|�ab,|����H^;<���C ���^?���q�`}+�����Ն�<�k:��������[�s=�<��G��q�{ �O�'���q���C%�]2��~�$��E��\#JBP�{y�c*���,�Q�!���0��������3]v�Ex2�n~�A[�t�����d���S���=y�(�# �5����Td���%�1�x;>�x��
���5&���5p9�z%���p�$�G�T��X.���
���t����qe1Ύ��m���$�2`GF�u����i���6�@vs�����J�Ɏ��:I(�6�J!$���P���]��0X�.�=7w�suɐ���(����kE@�2��(`Pץa�&9y3�:���v�>�T&J�Qͺ���Z1�g38�>����q	%u�Ƞ�u�"8��r�`��kV�W����v"� |���؇c�ϩ��X�v9�/|\^)�t#&ã�_���L���V!"�Q�� {�΀L�i��H��)"v]/h���q/��;�����������Xľ�׆_�}��S�bn�r jƟ7��cY� ��y~2��>U�T���*���&Zaa�+릁���m5v4���}��[�e��_��B�+��$`:I˰q6�n�1D:��R)2�����q�Ym��
S�ؽ�,�R3��ˉ͙Kw�}�[��o��q��<��H�i�-�kh��]��/�'sZd��W��� ���� �p!c�v�*F٭`CNka�.��?����a*Ix��_�ȋ��d0s�/#3:E���C%PO�{|ބ6���n���bRnR��6�8T͘O��L�u�l��������#.:F��U^3�A�i����F�H�{�y�S�%��� �R�S�qRү�7P;��������W�����d�;i�B�-G"B�˞M?>o�l̵y�Tiy˄pZ)E0�w@y�!��ր�|�.�+�f?��}w�I�̱�<�,7���p�¹�8���vo+�zN9K6�t��r�&�	��sڙ���p�[��)VF�cM�o{�%S]k�#s�j�)�5�� ��[&Rn�_	��X��(��h��An�״��?J������ޝEϺ�*N0�:O�K�'E��ㆅC���$͵�:P�7I3tD<z���q�0 ��Y!����blܔW�{]�j[;�A/�.������"s��g�>ӌ �|���j �堜;w��oOLZ�� ��ÑICrIuuj��-����V
~q�m��jy+��%>ο�y1�\�d�٩9�7R񯺹0>�G�9�c8�̖:�K �ay��p<����$�c�Ч�� ���xw�YA�"��a��V�e�=��K6Q6��^׈<?p7;��׹,J�D,��Ļ��[�":<���f�)J�cs���v����~�P�*�iI�m��);�A.�(*�����?O�3���T�	P�ӝz3w�&��~���?*��wI����I�/�K� k�4���P�0���YdQ*�{5�+���(~�#6�2���e���Α^��zp4#������ZZ���m���������@X��l	��򗠅ݜ*!f�Z�:�,�mI� �EZI}K:��B�ݻ	��� ����n ��V���^x�I��J�(�+eXշ�f�	�N��[]g�O"��'T(TU�;S��P>��W�DZח���/��觳t��GQ��Jk<����KLX��S|�q��th	}'L������Ia)��:!]�
���X�����-�����29��Sf�(�C|_nk9�`�x6���6�j�ń?<�����kldަ_P89���;F�8�-_BgM���� ����^ng^6.|��������O F	~�1�]�e�׾[A=�s�.DRd�FB�2u�P�T��E�_��X�M�\�=(��~�3+9����-��(hd^ŋo7��xЗ(�_=�Hf>�Ҹ�,z镗h���L��{�U7NxN��Q�qdK:���`�I���}_2i����=[�5}�2h3�	ΩiR��B�k�k�o.߸+܌���Û�w�_Kc�$m^^��2�r�b��&��L,�� �*�>Kr�1����{���dd��8����^��I{n��p"�Y��X�}gzby�l86�-mwf�(=��ޫ���B�6����W6Z��˒��#� ?���0*�t�X�dô\���ۺ��A��~�.���+p ��{���.]��$a���Y]��3��s�_A\>�nL%xݘ�p!���>�f���/�j)l���085$�2�?lC:^t��;�IsP ����!����/���0v�d"e�º�u)
6tg��i$w����;���}�6L��#�#�5�(��ƲPe��4Ctm�}�k�%��?l
N
���5�����R7ۃf�����랪���Q����>=A��;?��!}Ӽ{k{G�Fs��T�A~�{��Qˀ@��?j贩�$/�_����%8�B�ַ����[�"l�a�ʅ���W`��j}#�K��W���:p$��P��ܒ&�[j�������'PoB���т�e=��:u�@D�^���3�����#�H5^	M�h�Z���+ݜ/�фN��k��~\���}(�4�b��kT^��mi7��Q%O��n�ţy�}��/`ȿ� *���Ƽ�V��٦�T+<sCNT�͟+i.�܉�����h��n���� ��F�
^Bh��8#�	�}�>�	�p�<�L3t�A��Ё�
�%����j@J�E�%x� ��į��&�r���l~�2�8�%9m� c��F�����aA�Ka������jae@��_F�y�K7���'/��7�)�%Zr�I228�xg}lO|\��_�����j��&���� 5���巅�2x��+\�C灖'C�}a��n�z�w��^�M�8`*+Ky4��� G�<s���t��[+�C+�ᱍ�'�q�o�%���N�幎[�4�L�\΢�*`֑�;���?�g���bQ9<�6O��l["mҒ�t�z� ��3[�z�5�$�Ehzw�Ŗ*�#�,me|�MK�x�m[��ګ�Ǆ:#���y���< �^�dr��E�W����W�8*vl��5�"u���k)�ڕ%�t�K�t.��J��،��ֻ�Q$ ���l�M�[��n��x9N�Y�����fP��#x�T����h�ʧ�!�o�OC���g�6�=����3�k��N��f�Y_�p��꽭z�i�Lh^i�m�[��nJo�����ʏ�lO�.K�Gd�Mz~�!�t̵3"����������v�&s����=�`�;�(b�w���w6�a�X�.��1��Q�����udI��!r����G�#��\w,F~\̋���
�]�/~����͆��Z�8m�t�����~��<� �@:�>��� ��YW7���	�(\���(�)��t�[|�W53�-� �qb����s���ǕR[ֺ=G�Sd`�댛�=���s�b�.�e��y�e.p�bE~TT>���o�x{�z$����\���1 ��6�=�v�@�����vr٦�G���Q�K��\�����j�4,g�6:���*(���x�Rk�D����1�-��άP/�W�'��șO�6������r%��D2ߗM�E1�`�*qS��԰tl��x��}��:NܝB��	����)P��	f؄ƻ�b�3�QziЧ��e��5}����C
�!�+����Y�T��5��E��8�r�F�P���
=�'�d��]�t*��&V���h���u��:�G�4G��t��Ӂ�z5Σ�I�&���@X�5\�`������&��!��	��W_MP�\������c�u������0.��:v��0[Jw�������"����O���@��"i̡���>(���"��V�!`9[����ӊk{�DT����B_����u�7���l�� �������D�.v�ZZHF��X4i�}dU�\-���enM��h���?������7�+ª7�n�UN�����Ǝ�c���}�2Sh�!cť���y���1��Ԃi����k�~A����h��ڲ�3���|A�TL���,�Q��(����.�n���a��&�u�c��Δ���:�-��ߤS8t,ʊ�C�-<��b�(_A���5e�@ 3�=����AY�� ��C�(ҫ�xXLI�t4]���>v�={�t�^;g=΍�	�J��2��x��5���D� λ�K���8�j�(���d���=�� �}��Ya��׀�!���aNN$x��b��]
�i�r�h����~��v���
S*g���Q��D(v)�Z��$���,r�AU���2�
����t�(���#����A�����=!*}�$��	�����R�?��`����g�$�yĈq84���L��g1��R�J.f�9`�
3]u�?�KF���vM��S��\�sqS:1��P��/�+��P?��Sb�0ig��h�L��^c�6T��z-��2$K6��w,��^��%wҥdr�ئ������IDd����u�)#�} '��@[lh)���$�{�.����:�mA�8n��H5I8F�3i��%�ҩ���?���'�BX�Tm���[�]�F+y��C�)�|Z�^��L���D�6rI�.3Ol���3(����I�����%o�d��Y�\����DD¦5�}}%���Q[�L�R���N�(��zmx[\&�
�d�N-���m �w7(�-�$r��mJDm�J�;��(����wѕT��b��Tn��ڒn���3=��eȀ����p� ��۵��˰��~�Â~��ؐܬpAM�F���M��o-?V�if�Y�Ͳ�i*Z� 6����]�}��%f��a����޽�T����5*��Oc4����ʕ�sjH~ZgtJlַ���rj�r�uzLb|64$4#YL,�[ڒ�ia3�`ՠ2߬��T���p,��5��7��p���q�Aj�LG۫�U-W�͋z�fȢ ǵO*���w\4��Oz��W^�z͝���,��JÂ@�����k������/�I"	Ki�����u�����~�75�e��ux�7�Ç-��B�����0+_�{�i>��Ţ���� =W+'�l�)M~[��v���\�������え�&n���_��?׌{�t ������Ӊ�������=��͜=����4O��^�/�89�1J��z��I'����o"�H��Ѯ'e@�Fr��=o���I��-���5�îx;����]a`ޜC����x[������9ޥ�Th�%��ܗ� T�%���wG�۱�L0�ǲ�L�҅L�'���i����r�,������aK�����K�f`[]�(���P�hh�H��[0�vv�D"e�����^§p��C�
�r��@�S�5��6�)�S֔;���j���A���F���5�@s+#s1T�u x�Dq�{@��MTO'�zc4�i�Ss�~�uIV��j<ȿ'�����?�X�E}�Q�d���X\g ����a����<:�8�$}(IE���C-_��m߳C�N����^��
8K�W��T_~��w ����C1�0d"M�߮b=e<�c�w�ɸ=�V��ĭ�,�V��4��!}t�s�3��^r�\��km��Wyn�<)D.�%��;W�"O��?��+��s����/+��y�^�OK�p�Bo�xŗŀ
����L��� H�� x�s+B���U�	Ң��5���ѫt�x�^'��ӽ�T���j�>��z%N�v�'ft@E/r���.<5t���U����A���1�0d���L�I�+Ma2$7',�%/�YMG���a��/.���	��\��v�3Z����B�b9�Ç��3��5����i~z��SM��ؐ�\f��<G�$a�R8��fj��U��$̗��	�7��8�z��V�Z�l<��9W�'��D4���'�+���=f������+�No$���~rU�Uq����lk2����γ�u4a9K��_�a͕���S��E�U��[��&�E�B<�Ǖ�)=�CG���_��$�'D��P�*)�z�.���?�n�n_��JAq����|��Ŵh�W���x�qkBA�".Qm��< y�q�&��[B�/�K2��Q��F����ޙs�C%|�N��D	R�]��Ӳ��5�^QR��nT�_�)z8$�	�g�v���#)@4ˠ��!�7�$��%|����W�>:�k1��O����fQ��F�t�N�:�*�H�=>���(Cs�� {�"�dem�l�9�Ԇ/�5� ���A6ٯ�mP"#0р��C�r�/�Ia�M)����xW��.GGA�583x�Gy}�T�'\Ć����$��0����\5��U��v�����e��(؞7�I93D��)�g�K\[c��b
Ca�����.N���0�Z�~ߟq���a`M~5n�~4�G����:]��W͘��6~�f2�)~�Ⱍ'D���o�4t�MR�����j_3=�+����g̻W{ �ķ�����M"�~zm$�{ʋCR�� `��^eT�-A��ɣ����g�R�P�j�fF�Y	L����g/�WŢa{�nϟMOh<_aIn!"^~�Y���o6�M���%�L��+�Sd�~�$gZ�M�ap�o��KlC̓��49y%��`�K4i�+5�A��5����U��(�X�,����Vp��ʓ�ľM��6�@
�+{�$�L4J5o.C�1������8�n����fV�$ު�
6[$�I7�3�
���K���tM��^;��HVȤުvF��]��P9��׉��Z�0)m�L���<cAC��C\��ӰNA�ӂ��e���0�A����-����vH�2px���o_�H5T�����������ȣ���.���U'�o۸6#a�H#�:��U� ���}�̞ᤎ�X����R�#�FͰ��~L��������?��r	���W�v����X���`2x�\@�g�XE��u1��;��A�w�������jg/_�(���eL���-͛~�+3�^ ~�z3?�I�.�+�|ֺa}�n���H�'���Z�!Z=�8�p���l#�˙i�z8�j�jٚ�4�F}�V�I&o�R��SCQ��+�$����H�Y���	���e� L�����}�큇�ͰM�X�-Դ��(�*�>r���L?*{� v�MS8�Uq�\x���ަ�Z1��';�ӗeU�n9p��5���}?/*	ӟJ]�n%�uk�L�3ť��݇��3��U�J������;L��Cv>Dʒ۫�,m�Sl7c���|��f��)��n��3	c���?�H�pA}�Pݩ�Jl�*1��͎����7�nѻ��e�=����\�͙YStZ}��Uڰa�,��ΰ1/�.�^�Dx�-�@�z},��
8=J��;F�e�kSkfNCd����!��eb�l��[�i��B/QfB�䡜�s��|F��?9�"-��)jFi��mjmkS���y�����~�
oX꜍e��Ctҩ�7ӡ�?.�L���Y��>&�?gg�w�o��*iX9f$t���J�\���S.�;LH��!�rR���]��^�2�����&&�>�sz����`�{*���QK q.m����\�Q��� ���3:�����N�-�5 nI�V>F��J=��~L�]�u~�EQ��ڈr�>\�t�����
-��Iv�f���9�r��LT8yJҏ�K�7����ʇ1+T�S��pGu���&�s�2����d����I��p��e�ie&bY������T^0��yJ������`�DDN�S�#Ր���?�E��uʸ�y
��y`��fۑ�E��4���뢼6�����#Z�GB����K�
�;���	��\\��� D��*GM�s��:������m�{�4�B�kn�!Qz�J`C�h��6�w�D\ZZ��	��tO`���3-�����a�}�� R%�M�G�n�<�:p�#���U[������O�ǻ���`XG�k����h�������J����o�nHO-:����G#������t��Ի����$���k���XbAȓc�L)��;w�k�m�wq̵X*�+�b�A\��&�˄q0��}p�/�	o�|<[���gH�R퀕i*z��Xb.CQ;����E��5�˂�bw��"���I`v8�X�io-��l��q�,^:����G����{�c 7 �}�V~����UY�#!�j�I�L�	�Rw_%��0�Q)UK�:gW����H?�4M�e��II:�<�'�/րQ�V2�N\��r����P��Yֲ<��N���F������ϟ+Ax���
7	%�ʨ�1JBF@&�_��zA�y�y��������z����Uk��Jְ�k�Z�Hk��j)5=��/ΑN��`����nΣY�T�y��/\����gTS�LwC�U�~'����f�E��R�ꕢ����Kr�҄��eeTR���*'?��g��'Op�5oҠ�R��c �;Y`�j83��b}�|��� �<�K�oɺ*��]l��f���{v�m�m�$���T	ݿ�7�P8��k�:�J"�8;�?�G/늌&_��q��~7�A�)9�񬗻��
E��"����D���AS�` E|)�I����*���N�3�|Y�>�k�V�6� m�=�^��K >����A�V���[���9[.z϶}=*�xo&�Ԯp�^^��#U�5�ǆgG��9���~�B]����`�^����3n��Je�>~t�~aNB+���P��5Q��Q��kN�@����Ti�����c��3����ƨ'e��U7Fik���%�a��>޴b�	�iy�W�?E��	|ޡ	��4�O�?� r"K��Xs�W�{�`��s��8��o/{�2.����Laێ�=�	�K���^SC�9��#G���=M�痃
�6N.��3hR?r�V�Q���}���,~��nTk¥��6��R�OI+7�3H�#f#^%E ��Vҕ�\.J���z�A؈�(<��K?�ꄻ@�[e��:{��1���8��n��eΨ������Z��i�.�Ā�I��b��qfZ;���7ir��0�����y�g�Ib��S����&�ۿR�\%�&���9��)����+�6k}��l��oǘ������{6���������j�x�hv�}����T�k� uӬ��W��2LÎc*�L*��^�Zwh��ӓi����L��y�ڞX	�[1;U���g^q�7决��z�/_�>���3+M%�q�(*��Y�+�a<V}��g�>x���Z�����V_R��B)g΀���4�R܎.S�N)�h����3�`��~n	35L�ٳ��yvO��d��$��|�H�}�Þ�hiL3��_�I4��W�e���F!�,�K��?�w{ۀ�={��޷n2u�x�r`���7�&�t��>Sa�_:���R ��&CI(K��M����M��,����Fހ8������=��2ԏ>{��l�����#������2��#�P�Ӓ1*�P ����00���b���G��4#|�K��h��x�<�ـ���qR��n��dҴ�;�%��f)����LiK/�?CT���(��[=Г���8)�����(�&�*��X�k����ا�z\3Ïѓ�;�{�y�W��� ���b4t����:J�<�Z'S�_!�%�� ���&)M�	��c��U�CY���7���5I��$�JE�����j��EP���l$�"�&�a�-`��F<)��>+������-��;��
�	��&�Q޶�ڋ��N��a�3�x��� �[����b�����R���L�U�X%kgE�W�#Q��iZ�f���8x����\?�H�X�:�g�k
�n��Q�c����݌Y=�/A���\2��P"G3�ul�u��pc���=�$Q3�������[m�~.E�'B5����Gn1��Pn�l@��2
cP:)]<s8����=<�jv�=��_6?B�=(R	��ԙG5 I�H� �-ܩ�+�%�� A���<�����
�1���H�>��Rf��\���>�r��;U�����7"=f	M�����Ţ�w�5�ڣŃ+�tz��ґ3P;�Δ2��,��:�8K�3,P�I0�h�d �ص(�k�uQ,0� t\���4��ǶD`�Tw��_h�����I���fn�`=	S��qW�W$I�� ���s*{Cd����i���ʿ��"�3k��y�	�>YX�C�7��J⣵�����q��d!��ko���p_B)�k�3�$D�	ײ����	a�q�' ��������5����0m��܀Ӈ�x�n���=~�ߝ�>�$�O��)^<x!iw������O����y�-1�>��W�R_�������dU[Y�,4��ߓS�a��C�Jj�{B��f�����(_��3����R:���OCR�Y)D��X]�R~�j���
U��M��n��s�.r�d�4��XҩcN���^k�)�
��!�C���)u&�p*�V�i� =;�y���Wޒ K-AƳ���]j�E�iގl��b
�jX=:�_���߀�k"�kEL� rb�V��-M��&^�+�ac�����=�%�TŠk0>L��Enoig ULh7� �)��=����M/%+��9q��m`ҩ
�=UE��{<�2Ϳୢi5��?�k1� ˚_�?c~l��5��^0��H�.�Y�of��Њ	'gƠ|X�{���S��w-	���Ntq~�P�����	���?r�#����.\�������ldoT!������.9S�P���a_v�lo]�|�H�MH��#ہbbP���32�|w)qotM*s�h�lẄ�=�x��'v�ysgC�Y2ׁ�3�D�sCp���䮴�(Ո�Q6�bt��ǃ%�J	u �S�d�_�yW�)��+���}9��Y��c���zSc��ﰊJ(�q�<9Qq��/�g=
�E��$K;g�8��MLŋ����7L3[�O�{������M��Tq��	��C���,$��{���b�=��!ƙ�R��9�M��:=H1�l�A�}�ZF�]Q�`����[FL����w�#l��#)�k�^�s�L'�C.�<.:5y7���Y�r�dlTa��<��}c�6 <����.�E�X������o��v@j�O۶7ʵ��0_�8����qƎ=m���ASޚX��L�LɤY���!�3�-��Wx��g+�5���9.�*@��@x�`z&�C�{����A���\�B6Z��P���/��yÿ��ɰ��z����g��r}�/����"��}�C[�0����́V(�h�ߧ݈z�)�o�1���c,�X˛tE��8�^z}���:�G��p����A~����vb���y0�2���x�ۤ��uq��/�ʌɻ[ŵ&�b�����Ϡkr�T�8���l�!'0��dg�u ���m�3"Lt4���*�q���$QՏ���t�5�K�Av}߅a��B�͉�7�
	#x�O���u��f3��+�hm�W�1HQ� <� �b�;�㏷C�,��fھ�/	�����Q��[���΋��uG_fu(�$�[����Kõ-] y
'�ڈh��
-��uJ��j�=|�b�LA��>�?���=��zZc,�S��끺�=�ݤ���K
M�}�_��R3���w�.;�=���{�ڽ���\t�ΐ�Y��V�T�!)�{i�����[�b������Ț���
������Q��]&�Gǁ&W�+���1_��2�o����\�Lb��2��ǝ^=I���%Bf��k�,U�H�_p��~s�4���eJF�t�ZP7�2�`:�0��{]��%5�^3_�;m���ID���M2�#v���P|��پ�C^�`@����1̐鷗�}1�̀g-7�����1'�mrDHZJ�S�����<�u����1�0HH+�S��B�$�n�	�9�$$��P|�T��a��$����JB���-K9�s� �6�K���{�
I?u�cT�h��*���Kr��ڊѥ~�����*�~�LT襧���p��T~�E_�s�)հ��hY����i2X�s6��!��<~d�3!��Ub�4ic�Z��`�M�v*��TX�4@�;+��jN���j9��nFP�� ���q��U�t�iZ;mڶ�1q�9�eay��R-���eǖf�7h�RsT1��΄h�� 82�L]�X!�jL;Xw>���j>;��{��l��(�f���-V��W�x�/���^�����!�	�&��m}�j<�d�^B������aeWe�H5��^>G��:�}�WD���@�xI{�w�����o1�8Jpe�O�w�Ҙ��}AWyTq��6wCb8w���n�y�����,qF>�<����{<�8�=�(�fh�A]R�\h�� ���|a�����,�ȴ03r�l�6f�#�K�la���Z�
u+r���g~�q�YQ��H���3���w�r�y���U�~��;QD�@P�z�lL�� �v�'��-5�A��R��N�, 1Ҹ�Q��;�PL��ϵ�#�D��sR�ˬ�IFC8�?�5�^���H���2.��.��������m	��{F��-�:i��W[������0�Ux�=�wTD��۹��2����%��J��!��1�vˇ(�_M-t�x���CrW��� d�'eL�d"��Cq4�7����T��n�u_J٘��xPpm ���m�OGx�E��=����X��X��:�\!�2�
gC�q��gO�ȑ]&䍍;
�����Ժzg`�MEl��<��4����)�A���V|�[8O�':�ʪ'q����������*�mY�)j�I�]����>q O��w�2	E<Jy��[��׿Ϛ~��R]�[�7ΨfPu��CψQx�J���ن�����XҞ�~K�r��9�áLd\�E�bXKƇ������I�C��f��'�O�e&�׸��d��~ߡ	���?Á]R�<�����R����|=��N����M7���K�+���R�]]�G&kY�L�D��h$��ً��ea�I�D���o�� i=g�/�8q�7yM-Y-X�ߨS�S�+�n(��՚��I%���N���#~Z3{^<�����%�O<���F�����5
E� 	M�?�lOA�\x�qT҇��B��6����Nl��}��q�#��
��^�j�O6�J6EA�J�����$�,f���H�K'<@�x��,��-�J[�#&)lϿ��x�������,���~V���}�-��՝W�Ѷ���j"YX��)�
IaД�GQW0�MІ��<�1�je�'��B�%�AVF��Mc�7O�m *@�JȲ�@�x�Ix4ǈz;K >e�2do�b���j?�$���ve*�l(_���$�Tt(�@G�&�P�&o��w��X:9k/�z��M�x!>��Ĝa�|f�DO�j��b�?=����q�̒x��a����� NS	���$�vG��l��
z��yi��:m�������fo'��F @��
	{a�RN��0����:x�&����|�u?��\��%٘p��Җ`��|�j������d9��SSs��b�N�Mw�(�^u�G�B�+ �3���ڌ8AK~�*����i$"��Z�u9wh���Q��;aO;��t���z+�ȍ�_SI�`��Χ�d���oND�̔d�$_Խ"��bqN��d2޷�_�۱<����1Ee���X���m�f�Bɉ�f��8d{�%��c�ķb��H�yp���sJ�SZY4���C�b�Sy&�&x�<���o�F��K�1۱JT�'m�4ۉ1Хk$�TL.�i��m:�q�X2���_�g�r�I��H���[�T���Ӏ���jF*l�!N#�5ގ��u�$�J��qt"�����&6�RIt��Vな��N��{�D^��q�:Co��S>�j���ɧ�^8c���8
_ޢ0!#�$(u���aL����xumC$��g��e�h��xXK��J�=�-g��A[�5��8�� �?�=�t�fb5�y���JevUF����ȥwc_�����_��w�R6�5)�a�Qu�O��gF:)���@:z�9=���4��6t���Xt)dDy)���d�6X?���s�sI|OZ�@��rym�1
Z�۽k���������q����B��舔�RS.X\|���O�9Vʴ�y\���|�Fd�!�>I�0���R8��CPCC�O��މ �؄r��*�'����0�%�F9�����bK�t�"x�)�hc����̩N<Y -_ݷխ��X����C(��o`���䀱cp���1v�h�,m�,���$��@S+ǡR�I�Q�"�6�?���$�J�J
���C�-�� �!�q5�[_��
�@���.	�e�	�n�k�� �]�����4]��^�T�C����Dk��3+_� �ݗ�5�3�;��,z�,�� _�\k�$�������;\��p���w�[@�7X.�_t��:#��;g�U�{t8�X����q�����H.��.����['��7�CC��d���?�Tp����@�r,�y��O2LD�̲[ܽ�FV�C��tZZ6XB>Ib+��9��2x�lhr����:�Kc��ze��{3�:{�l=-��.�eV[4���0�R��i���i���+ڢ`�_H�@�)M�E죴���:���ߣ�Na���*zr=T�X{ƫ�~����c}W\�F9�6�ʑ	�$�;���iN��,�܃Y���P�G�!@3?!���9�G��>!w��7#�>�1|�t�`<y"����Z�����o]�<�w����������T�(�z��'��5�ut1��$�x��0�v^!B@uţ��1�y	��D�N� Le�~=�zc���Y������E
=`�x	�����Ra�o�RF��������T���1Di�6d��K�����yg��J���F���	��]��uM����lwϲ�HKk$h�cmRE��o�	;VT�Ҭugy���Q����p�֑B�h��h�Q��y��p���Z�=���k���q�30�E;��&.i���3��*b����~t�ٜ����`c2��H�Q��-�# �%a��ˢġ��S����
���`��P��䐖�3AE��O�ܓbuA�����ޥ) �F��	���Q���qA-YF�yc;D�U|�E�_�sq�Y���L?��m��A��Z�>�[��9f<O���i����r�t�� 5�{2�B?�`!y�`�~��t�\m��JpK[�� ��X7�5wH�6� �>X)8�����L̑8O�zl�u�ķ�\�J:n��,�}A��T���k����_LT ]!v�oo��[[C��u�6�\�����Z��hX�zdgpv�=���\,��q�ۼkB�]y8j 6�������1�(�D���0VP��5!F�2C��Ǎ��K�]���<S�*^�H��}߶����Ԇ	 3���P{��L��Ib�G��]C�}5�u����%�^��t&�>����.��_b�����b��\�>���d��Cɴ���`ΪGKۭ!�~����ط�H�����&��L�y-�.E>�]��.����]�=\KV�o!�~�؁	V<�A����t ֳn�������6��ⳛ�y�MaJh�I��k�v�0�)���C$�|U�8���\���G�8&�,�K�q��n���g:5T�@	�4��-�� �/�?S��y��	�c�� ���g�kuؒA�@��Cנa���_�t��dH�d�2D�K���ʗf/i���,��;~�{��?>?�oZ9��ǋ}�'7{~��&�7�#�e�����<7�������%x�G���ˬ�i�s���<K�6�Gv���WLRi�s����r��A�^�|sl� 	E*׳.��V7�M��Ou�퇮6��x��^"���c#P�R���T�K�¼'���n����_ծ{A��2�6��9z�;/�����d���.�\=S�<��5����	�m�<}���Učn�ٔG�O%�yr�<D��rO~xD��5��R��Q��PN[�2�?���!��}/�U�~}�C꣹V���RP4ב���(�B�� �P۬>�h����ʇw�	�^'\=ٸ���23��A�<� �0yA(�w3�(��$���]� ��@ǔ��G�@�Zhh�`Vww��#��	��1aQˌO��|���ԓ�w�����	�9��Yl�~j�c"��={�.òeoX/w�fg�ڃ��Ցh-�|"�9R���Z7��(��,M�f,\ Z��� �2��B9R@<�@2EMn8�w� �f�r��#�qu���k2�r�M5�3�Zq�`��߉�2��.��h��:[�lJ��S�\|�]ߺn�$�Mȶ���c#IiNQ�A�	Sua���a��?�>�6+
��N�t�;�|���f�����r�T2����=������ׄ���w�A�@�r�d�/���[!ΚK�؁;W���8 �w q�
Hj��E�w6����8[���_�b#)?�P��2����edE8cw�?\@X��B�V�K�a��ظ_ײ�X��C8�Fq��6�J����]�qP�tD�@%�F^6IZ��﷚Y�`i@n��f!!e�g���H�a��(A���d9*P��\Si���˽L�px�l���ӔToضb�3�=�w*��l��s����44�v������܉o^x�xx"x͗���ՙ9_ڎ�Z������i�I@��2�UQԚ6�2�;�Z1.���5�v�z�ͪ��lS'���&���>c�w��Gئ�<M,7$T��w_����"HS�~���ƙ�s�؜���	d�v�]Ĕ����Gv�J���ď�.9�� �I���qqϨ$�����R>ƣϒXQ����K��-��]� �TL�Wr���6� `��r�"F��YUO�Rr�&����-����Kd��
	��+}z����a�ỢӉ?�̈́�2���d�c��n�R�S1`���lP�B�Yx �EgSz:�L3�KGd�U��5�l2|k�Aj�q��`�g��A}�4wp:@Y��I	:�A@��js��nL�1���q��������#)*��isYv!����ԇ=w�+M� �^�V¿Ǌ���c8����&S@�R҉k���v��#E��q�n��%c�7s.��b-�V�K@5�H=&����+3J��4�%�#��-���KdV[����t]q`���d��w��$sֹ��r�a��-�?;��NO��iZa'�^.Y,lѷaj.�w�"�z� �5�!�g�`�3���яo)��ufg̶��K���4�C��� ��[��	a��K�̫�N?�/
��v,�Q���|�[p�� ��M���f�4ĎP��輖�}�0,������~��B]�rM����Y���T�y�[����x�O�!7d�̭�9׌�l��E���+�1����6Bs����%b$	[��FuL��DVqY�V͵QT1��-W�p(�-7����;�PopN�>�ӾK5㧡�#��8���[`$+�lX�2AX�`�ҽ�
%-���3B;�V�9#�l�Ő�2�A6 #W�J��ն��&ח�'qz��y��֜DD��9w�5x׮fΖ	���2VW<�FPYRv��cRr��T#����߳��I��Y#�L��z2�` �HF�7N�DT����	EoX��ོFO��@��9G̑���]u��~�8%X*Mp
 ����k�/'^DW��H>�=߉�6��.-�X�
>�t�_{X⛞��A���N�S��.0�j���N[t?4�D���q��L3������	��7d��/��7:�HJ�4���O�T7V�ۉ��7�D��'�k�+T���A_��9�lP,@��?�,�J$�	��s�cѐ��Ko+�&��JHq;Ɯ{�s莆jC��<�C#ż���t���m*9��� �G�+�L�$��Q8�]d4RrR}�A.�`�C���v����0,w�����_���8Y���\]z>-��Ya�`�*,mw�����4��ވ�C�����z�~u�$¾<}ß�וn���I;_��R��xaS�����[�� �Y��p۶�I�J^}u56���,�x���*ل*Vw�Y'oh�Yzd��</l��ю�K�-��y7UO�,!���(�L���49퇬X�9)��\O� 1r����ި�P_�ߘ����38?��0�I�� ���3~(�bf��"MGei���@�r
Xu�g7���7�E�~����ӿu`��=@[5��xg�����P�qV�!t���*6Qجr:R�by��(�{��g���Z�O\n���s��~��x3:�0���5���d�:��=��@c�1�$;�gV����W*ۖ��
�;���b&����M�2��ḎP:���(B���&y�b3��}�ג$=��/&�pa��2��/kƔ$���\!������)1��<��7,,���Hi�>n�}��� h����25��g-`�0�B��0� ǭ�h\����[ח�o�$[9LZ4�IR:{���C ����S��޺/}�{J#Î��|'~�g4���܁��5�D��5.�/��7�) ��-���kt�m<CTn�o�׮�oqsK.���L�	V�ͷ
}C "@ ����0�\F.P���M+U�T�Z@���p�9�_�cR3��� n��M��"��G��37v�^MU�Z &�`��=/�K�/���I2ĉ�%�H&��A��4�W��ѱ�ۿoJI��y�����\i �`��:?�z�Zu�ʩE%�ZwJ�8,5z��GB�/"G}������:�)�bq|�+v|R�;�F�kb2�MXbw�Lx��25 �����1w�}�)C1�oE/��Q���=|�kݱrCE�!��I�G�J&�샅�#�0�w	�\J���ңo��/F*�l���&GP��)�Q�QtG%
,�݋�W��n�<��Me"m5���pɪPE�v"��P�1k�T� �
�a�+��Ot�bٻ<��m���S�B/��J�*�&���-���S��2b��P|�M1��[^�3X��#��>WDh�E�>W�x�WQ��ݯ�\�=&p��~9V=��+��ۼ�!v��BԚ��rÒןbt�{�@�D��Ĉ�ȣ�Am��v���%�쵕L#Y��t��ra�h� �>�-���F��\�TY>�S�����u|F0h��M���ߤ���a>���my'��16I� ��@����[%%7�Tl�Z�ҷ�PQo$���ŋ��jdmm*�?��]{��%�RV�8��}*�]���7����%Ve��#1I&@T��A�)�R�M8=ū����H�rYȨ�Еtl	�Ǯ$w�p0C	0�t�Bv�A&5%\$I�@w)��i�x���EHS���,@ßv�oeq��CG���r�uL�G��/��%��
���u��gC���PIsE���'� ��^���M����cZC���L�r�[����琥.����2�]
%��MY����5�c&��bH,3X�@���L�9lV����j�.
�J�G�[]T�Ѿ�|���T�U��OP�↩��M�]-@����`ڿ��d�*�(ݜ��4M�8��b @&(ؐ|�c��ɀ��S�����(�i#_�Ty���)M�|��M��o�
k40����=��~�!����-h5c@������ d�G������!�?S�Sc�ƴ��r�C��NJg%��!����2~݃w~�3���L{�ݲ� ��(���k%~���'d��li!��G���ϱ��*s���o�������t�� ���ͤ���G��d�	��Q�� �M�x�e�ɰk��k��� �gd&��e��G|��˷ѣ0�1�������H���Q�����<���\2�y57��m"D4a�뒹�����wXH�_u3?i6I�:�@r��Z� �*������ ��o�:'�^��䱦��??IY��)�6^�M=�rփ�}���I�����|J�8���!>�N�À���f�rE�V4' 
E�u�+��f���Q���,����_�[ð'5E��*J�E����� �)�!���!S���f"�ՠ�,��R���cʃ:[5@;X>c���ʽX{�iÖ3��z4���9�˜�n��Q�X;�����ݵ���_���K��*�1a������^��Q�ۆ20_��-@�5%s�x8tMt�D�:�2���*P��bPZ�Fո��ӈ2�3-�`Y��� �j��B�a0e�JЯJi��1?~����=��}!��z��P� F��a�bڌa�Q��C{�Lӻ�;�B'Y_��+6������H4� <��3��`�t
���M@u���.�U6�63,�|�/ ����]<�ܟ����K�t�,:]�ᄂ�����ἅ��&�Zlb�gݷ�<	��N7n|�Td>!�M��>�rpD�"Ţ,O��_Q����ݾ��㼆`C4`�~Q^�3�����Q��K86���S������`����6�+�X1�?�����aI��$��Y��{�w��������RYx�N����R(��|����L��k��a١x�_��

���$�/=Ro�ԁuc(�7f����YNd8C�ƕ3?�����uow�8qܪ/���.���=�	3���������:w�d-�[u�G��b��xO� o�ܛ���-�����1W�9X�����erݡI�g�:L���fN��&݀��$v��!�g�0�a�dۋ�ƙ�|�0���?<	���b��R��-�%�-������Čs2�i	'ўx=VC�~Wa�ǵ_.��t͵�L5z! W	�6�N�V��:�،,���.��х��>Nkv����m�������Z�I�|7� ^FD{�Gϱ:�T|ܷd*����l����s���i��d8�f�&���
���;�W~G�	"8'�j-�(�M� �4��U6Up�UҎ&ɪ+����I��"�_�[�X� ����H��t���bF��f
��	�<x!�솃#{J�:�y�`�u�����'�ρ_y�C�8~bڬ2U��x�O�dn��,]����G0C��c�?6�&T.;�A9Kb��"v��6�_���qP�����'%��Xl�od@������Y�[v�&���[�N"�l�����Ԇv���>W塐��8֓�'��p�*�$PbY��<52�nu��6Blј:!�0l&܃~��4=m���6���6~�"]52Q���]�O���t�c�Ǳ��5�ݑ�$���oSV	iZ����GYR���g� �/��9����iu[�j������a������Y�:X��-:�O6��yI��;� l:UN�$����?��W3$�XR��G��!�y����T�X�۫������ ��5p������^������5��}4@��T��ߟ[�plT��.8v.������Y�J�G?����GQ�]_���R�#(FJ�4�OX�=��-T����IXF�2�l�L2#�Ii@�zx�ɢ�&(yVd�ڔ�ܽtѠ��$�*��U3�Y]0G��N?3Aϊe��V٥O�
�?��m ��OS���	�ߋzɯ���su�q�U��|U�h���� N���7���a�������8�:�2��)��{�=��nOi�&,t��y�b�q���@����a�t�:4s�6M��u�����T�	Q���n^!���g�2.C_�>�R�$�i��z ��Y��@tG��҅���'[a!mH������C}�g���֯�Y�&�����u	���w�z��HAO �pF�@8HPA�����&��������)X$HN應���J8�Q'�.�v�������de��H#��o_}~�Vq�%rTe�F���XZ��y�Y4��$��Y���������j+�;!ڊbv. ٺ`�v�B}m�G�v�������o����G%x��j��$ΣZز���^Ƥ	4z�:,.��U�6��Z�����&�D�86����V`����� �4A�$iK��rղ���I/��i��G�V��a���W�N�D}��ć��wǃDm4ɳ�gI~3U��ȊZ�$����!��,���۩9�H�ߪ���9�.���)Y�?�(Ǔ����Xƀ���}�N����-IO�KZ�a��}��W-c�җT��hx������T[�t۟nAg��^�3vk��n�.��=[�����`���k4V�-{�Ʀ&c�UPQ��'�3Wǭ��-)�*�͆����G�!�T���%;f+�b�պ%?:�뎣Ф�Ex��]!�n�j�]�\��kɤ;�iC�����J�ߩP�D}׮_Z�^��)�^6�����v�<_9^g~]Nj6j�m(R�(j@�Pc��6)�u�d�0���s�=b�S�������Gӹ�<q��#6�k��Q�S����`"#ڼ����u2=A#�i#d:ҝ���D���/��JY� ����B32 ���f6����� ��g�v7��=s��A?\�����l��L6z۩����ʔt��ֺW��n�=����b����1�:ca�\r2#�1R�覱���&��_`��ɳ�E�k�0?�B��K6�9OEExm�Ļ3x���.�&�צj�Y{�O7�2�N��W�蜵/�2�Rs�����±V1
nxeg��D��#^�;F&�a�%���.P��^'Ap73�
 � ��x���)D�\]��kO*����"��H�xa�j0����4ʸ�D*"�G:qֿw��1I���f�ƺS�C��5�S,)1Y�/�ն�~&d�}���J4�����x��眙�_8L������V�%qΨ��%=��.�s9{i�3�_�����~ۀ�Rv$�-���cxh��G���� ?���V��J�������ːE �4��=c��a)�1<��"��a>� �Vbl��A:�mH����D����'b]�ߣ�f��8�|�?[E���E,}@�0�df�?�[)^�\i2QJ��U�*��������"�o��YȭYf���y5zu4T���]�Q��jl�x",̊V��:Sc�ֽ@�ͪs]2n���b�>8Y���ﻦ���i���QC64,@�5X/2��=%�㹷�T0���忁i�ѥ��ȠM�l4�D��Py��+�yt����D��d(�4�Ь�#������9V�H��H�pZ���0nF-]]��"Q���K{�i��-�lL�)=��J9��`�䲠d�d��n5=�,ۅ\�+�?�߶Ծ%����D�2
��(q��~�ZaS6�Nreux<pz"�i���'v�+X@�V�`W�HAK&�"D���Y��e�4�F�k) m9����r�����Ǚ|���P�ʺ�~v��&A���ܶ_��^�O��vF8���2����%1�F����=�I�Kس�f|�.��[4A�+���W��_!��|v՞����|�tG,�\uf�f`��_�j+�l�C�=����l�h��?]�D���)�C�U�m @Ѯ&h��F�?5L0,jI�x����~���[�.��d�%V��*�P0˘�t����.�	���&{����׏��ӎ�d�l��G^�g `ѥߜR\M!s�;}2#^���ft�˃z*�������!�Q&��LmC*�o��F��Iu0&�@S8�!ɇw
�	ͦc��������� �43�Y��gN�q�Q��d��or��o����z�.�՚��4.��p����Ƕ��nG/_|�������q���{�,�B�CS8�9 p�0��4�尿�*��X�G�8'q]�X`CY�3JW����'s�oP�7���>��4���@�>���8��:�3�������;S뤋>�r��V6�]�}�(�G��/Ӡ���,�,�a�6�Jg'%��"&�ؐV�ўi� h`\O4��u��xmJ��J@����5��cD_�n�fc�@#xqGrv�y)�}K���L����)!�<���{nB�k�0�t�{��[� ��n%��h�*�r��>��n>�i�o����%�P�K0�;�T�RM�Aԛ��<�6)'J͇h�X N�1��y�]��匨��6v��ة<fK?�����;v������ݲ��(�0�̶ 4���D��\�f{n��`�6 ��ğ�a����p�r���'|Gp�LMA����_��N�	w�ar��.ϏprQ8�hC>�]�����K4V�>���˦JXiT�]�~��j�o���s2�$�w�Q<�ޱ�gAW.�t�#���F���z���� �S�����3��t����Q�~�A�1޺����o՝j����/�4�o�,�Q�X؇[b��n��de�p���9=�h��US�{�4��.sF��y�ܰW%J����z0�7��_�m�~�4b��VY�R�u�U�vhOSj�F%1[*7�yM�'��5?Ky�ȳ��`�%m����S ����ɝ�������{AIGe����:��(���}���+@��i���r�J�����x�t��O#[��kQn UX�Ӓ�\������d�Q��2�	��KʾM� ��)Mc�r�PB������d�m�3D��+��^Y�ˍ֘��@�^�RH�*]�S�T!/N�]{B��WcL0��T���RaU<v��vH�ۜ�J�ߕ>'_�L�?3�DG?[`#[�d�s�+��=d��6���Xj�	�.��(�A;��n�ML���݁B�M8*�������@t�
��m����|�i�W(xJ���5�y	�f+J����J��@� n�G'�?�5�V��!ׅZ�2ao�p^"�����_�d@��4���x"[��w'd�;>��y ���W��f���B���JF{�C]��!�#����g�?���M{�H:����ư�*�(��xq��b�2�JV!�d�����mS��4��W��<JB��&����^J�Mb3Q��n됒���ӧ7u�c�@-�E=URh\l���fe�.�l�@�U6����E3[]$e�:�ߑ��X�g�2�C�0C�y���8�D�X��OBZZ�q�~{�b��$X�I�> �+[ '�(���~�N���}�7/�v]`l���� �4�;��v�[�q�^��]���}[�	�|���7�T	V�==&�.:y����"J�F��(�v)E)V�x�'�@�Ȥ�-V��oFPf�M���a�L���������Қ����07�_�A�z(��������+S���:��l:((��,�;0�K �ĈOJXk�l�wl�|q.\K\H<�-	��'I�6��e���3N}��!:���[������t�K�=0�R!leӃ���,�i�ݒz>��ý'�{%l�c��$���e.S��Z�F\O�۞5,2���R��jH�X���6:Հ�V��c��	~��z���F2��,��H���r�� X}z�P����:�E�=t}{'Sf۰D�"��Zm<�Dt�������z�\	���Ȁ���$�WRB*d�fsN�)2����ς��_�I�:�d�cK�qŅK��� ���SQ��P=�нp���EYW��!�������uv���b�)ߩ9ƌ��W=���R�+,"��O�W�6�kO>X��$S���腲̄���fs�	7F����˾��EϬ�D�)	�cI�f�-�Ug)e�� ة��/�{^ѓ�"���Z(�)_{=Wͦ�cr῿��C�\P�8����{\Z�=	�-4Ml���M.�<��7@����o3�+L_�c�=g�F���0��q6S��	FR���Q�ÆpiIiru��R��e�s�KՂ�֭��m;.H���Xz�3��	���mn�竾=tg*2��޳��}�������e��'ω�h�?YkS�<���my	'�lp(k��1]��wC->�""��N�{dr�����s�?�V��^4�=�m-D#�G%r�uS$�j������g�Z~Юu��������瑃�+�LvOQ�u�4c�t�)\��Ǭ]�+��4��CU�,���UrZ�	��������$�m��,�T�NT\`KG[KGxT9φ��ߝ����ܞZ���9O�Ti�3=Y�i��}ԒA�?���L�[=L�����Z�ۥog3��(7\�P J�!;�[X���b{C�	��e@�%&��6 �-�#c3mU8r����8
����c�Xͥ���0i'v�Y߾�c�+K��/W�:���2��5�Ы�5�����ʿ_�\Jٴu��\�bC/��ڀ�sl�I'���똊��hHt���1"���!O�"����.���ڶ�I�����A��[tM�7�
�Pn��aDA�����]g��2��2kҼ��tK�N�<N&я��nH8�݈�/|�� �$B��ո"-��F3VI��sx��7��әߕ�4[��f��E������\��]e	���5�-���t��E~rmᄦ��~u���3
�n/�D�N^�C��咑W�&}{o�6�Jh��$G�~s��U�F��4E�·9_(�����*��Klk���-��堆�ucWՔ���A��^�Əi�=�_�{����f�N�����%��ƠX���YC��Ѹ�ͷ��ϣ�:_ZMG�>�.=�y�M��x^ޭ�(�z�p��7쐹��K�Z�p�v��"�d[��t^�J�_�5�Q2�C�>KH�+o)������;C'b,lW�[�בD.�a��� ,��'�?]s��k�hv�mE���0�I���0��90��kv��#n~��y�Ӆ�栶8	�?d��[�.pQ�OH��Yʌ�Kڳ���4 C�1��Q+C����q�%L�\`��~,���憅M����ܸ�	m���a�]������4���o��"�	Ƹ�k��:X�-�b��3�߁�`qڟu$ f�7W�0�ו�{,��kV�XR�C^�L��u!'6Cj���ƣRٺ��*YD �-J͓;�����t?n)s����C�_�H���� �`���wQn�2��>�Y�g��x�`/�Pd�vt��]L�W��^~w[n��� �B�)��WF��UE����0����He��G�9�㹋���"ҍ��(�L`G��"=ۀ��[�y�3U<X�0e����V��&�|13�PB;rdz�~9$P�C�Bq������d��NK���"��Wd����LWC�v�	��:��7=U
�x� h8����2�a�K�(��E)-��󥥯��ur� �[W��ǈm���"��������Z#�o"(�2r��|m�Vh��� ���j�N��x?r��d��0��\���@"��t�֡���"�3���ʈ�����27�7�phG���~�TaA���%3.{� Jzn&z �q���RP2b�.�%������i'Q�i+��nvc��/ww/ �j��u���oA��l�ޡL��A�u�E���T��+�@NV9o8��뤆����}9{�q�����&���_n�/5M1�����;Cӄ"2�۽E�{�,���Q��o�Z|����O��c��;�a�LÀ���r�f��)eJ�͇�W܉���fg�!G��p�br��d���/G|iڌ�$"��Y�u�Y��V���^�@�T����|���������[�� �V�]PGwѸl���`,��u����E��wo�����g�y���zb[�YDH�zg�����s�-�5�<�c�l���s`O8��)i�r萾w�݄�T�~��Mp� :CL~mM�J��k"*�ҐP�Nv}��2����m煪㥩t$B�g�$~��f��KI����MO��k=C���2m7]�)_�p�y A���r�~��xz�y��ȉE��V�
 �`J\j�]���e�M��h4H���sJMT��x���IE���A�����i[%>�C���?�mF�'c�����9����{E���=K��0���Cg��)I����]$`��y⨩�NAYg.�^���*��N��q�ɴ�Ǐ�v�0�B����q��z���#�l����4!�p|�d�|�}��)�
�s��f�G��  Y��,���NwO�t��Ep%��Ã,�HO�N�Q��*��VG�}��q���# �s�b��wzCd��*���EB�yXV����q_˖6�^;;XY'|:�6B�Y+t~�1R��q�<� �qΞZs��p�>Y���Mj}"a������|o�O8s)��o0��JU���.�[Ȝ֕|����$J;%�L�㽮Xvϡ88���O����<�ȣ�q�vJ����j��A���C9�:��	�dal���+:�q�ŧ��}�������Y�}(E�h8W�k�eI��x�$�ё~�ZɔBu?���䊶,�j-`��3�{N	-�.lsx�Ph�1 9$zx�-^XO�u[�EWH��G�"����M�7ˋl�Ce�$c�����<��%iAVo���CT����_������.6�V��[.�B�䏬�:���-�~��V��yL��A���3��t�_�K��m���Qk5��yϦ09��<�t��[�1{?����9�YƎ�1[9#,�����Ki�P�Avk�!)�y�C 騺���x�5���ͻ��M3BU}�%��!�R�J���`PA�T�iH��fy��L2s���rR�&�<��,�[��
�A��ʸ�t���uS��e���dř�7?%Q�_�|}�r34������􆗲
mW�A�J�����r:t��*�����z����:,M"������"C���k�����f�ô�m1��Q�����@���Q��~tWJ�nMG0o�U]�u3L ��^����o��5w������4#F�m�����ۺ3/�>/�2J���yn[���"���(�2��Ԗ#�`;���P�]&�kd���G��X�9BJr��'@�h��t/#��M�������۽�-�F�b�:��(f�.u���<x����q,KF�wE���V����-[,M�G�����.Ce��F�(
�J,ɏ�$xͩǑ@�q��Ȅ�Ԍ��/�����$GRw�:	����^,ٟ˖��b���LG�(�������vz��G�&$�����}!
W��4k.�L�o����M�f��������Ƅ��}�f���f�J,���
���Z��y.D@���v�l���}_E��j��{�OW�*H��L����3�<�5�ʺ(�H�Ɨ�k�~�M����m�vT�ɘ���Y�v�O��*������>gK}T��Ln�@s_�<��^�<7}z�V�I���+�jm���{�л��G`M��z��+^���Txp??&�>��w��A�:��@ c̩��U��0���cp8���D��Uo�&��2�tC0(΅'��%Y�*+��ت��q�]��6p:��&4����/�O�Q��EI�I�%��V�pB�9��:(�ɡP
Q�����b���F�����@�!�Us���B$Vi���r~���/� L�<�M�g5��5���H
��J��_��mW�('���YR�����QJCi�G���fo	:[_�aI��k����% @�������؀�ꮞ�r��eb�����*����MP+E��BG�]���N��Y �������f['�E�SHtGI�����}��R(�~�_U������:����9c+�����9@�_ң���*�r3i�=�mN�F��'�ې0&k�L�P�/�\M��W���/M����|׻��8uW[+I=O�	_R��y�>(����)f�5����Ғ��J�����7���@�D�sq@P�E$?�R��ӵM���
�
�E�ȵb�l��핕�.�� R�N��J�i���F��j�L0�R��D�V�Q��!��>f�5�,�}���A�A5���4e��:�ʘ �������v>��p���ϋ��d"��`8��W��i�-�
+Dvc�Qx�/�j۟��,�w�g���X��V1����&��avfx�0�ܴ��9������^r'��)\ۍ��9JO��=g$MH	qC�CZ�A����"ܚ+���ߏ�S$�U7Zӝk��,,�8�I_Sdp�˰@~����A�\7���L\ϸh�	�UK�>}��$�)>�%Ħ��n+T]~H��G�a��M�J��2M�����L����Яg�Sq��o��m6l$���ۈswVŀX�]����+��*��:�f��B��}��7�a[�)Q"�"���)+�#1�N�6�M������C���p
�Q���^ǓM<|E e���w{����*�e5�(���V�.��-|�2�BiKr�`v߱:��S�\����L,f�b`O�+L��#%��u���|b�[K��٪+#PITTs�O2�M�=��,[}�M�0>��[��|��饌U��I4;*%�����Ox�����W�O#�	ؑ뎎�I*���oZ�Z�D.3;�I� �����o�����nM��-���mC��<*8bE�f�n6�����fpI|l������͞�%�WT�T+���A'M�$�p���i�����mA`yL��%A$�5� ^��-�8�tw,��~�xH�T,ay���8%`�ܓ/��]���Ո���`w��� ���V�&�E�`��;4WX# *+aǇa��=[����:�������D���je>�m�c�3�ލ���T����Z,>��T�x�]����>���h29�ح����԰l��s�}���g�.r��]z����7ءP7[{b�Y�N��x^�' �?)��fF)�I�W\KѩK*jr�����dx!]����u�~������n�Ԃ1���۶�
���44�)S�����O+�{�{��7x�rF��"H�6�r
��,��V��<��G�U*��K:g�:O������L�[�T�R���"R�1��q�ڼ]�����Jᥒ�(@�֋v��X��i�xx��f3�ASrذU�Ë��Hn#lb�3Y��.�gvp����$Ւ���IJ݁�bA������6i�#��"�KpO�~�Öι��T��a����@K�h�k�����lh���+�!�z1@&�'�K^;[�p1R�q~ Q�O
:�I�ڪ�@6�WK��i�#;��</��*���v)M���*P��������;����.��t��h��Y0���r<���<�L+��%���X��yU��S���g*寱-����W3#�"�`�\lA�z���s�����k+G��N�rE+�߬S>ނU('����o�+V�!_���D_h�96'z����<UmJ�<<����5L_9}�F������	��9;��X"@�.0��6��q��S.��jX(�W�k"��a�.!+����J�AS���K�@5��c�3(����p����^�Y������l��S+�����I.+	�F
�qT�)��sB�Ҍ��7{Wi���5�w2�)�̫���a�cZ]l�́�o�;����r��reZds�b��A�+6�K��+��Xb-u�=%{q��|+9���ǊE�Q��|�=�s�Y�����`�ti)�N:��I�BU²2�� �読k��Z2���,K��`J`�b5PZPʜZ͚�~�k�p�����(ٙ���8��ܖ�|���szy��Ed$I��@��[��е6�C�W\����b�}+�../��0O�D�ȟ�q*.�L�Y��3��
iU�&uIz(hT���eQݺmu�gC�n����@$V���M����T+(�D�G��QäP�#EZwb"C�cX�5�^K*����e��xQ���V��˃��qCN|�hRa���@v�*��hlt��6��R���4�HE���o�me]��~�CPP/��T/���an�z��_�47A8����/��}�T`�?�������#��@�u��-�~f�h!��=�\��d���^��
)/N�X��;�Չ�:1)�2��0a�<3��b����ޠ��~d��Ue���A��I2�~�Z��ab=nD�d���8��� k�V�}WrX����k�g��]�C}��kjI�p���/]���sW�v%�.��%s�0��M�$���Oa#�>��/�Q�"�6<�b,,IC>��<C�ԭg�����΁��AF�7�� �M��������Bn�cC*�;P��5nW~J��>�R�n)�Ӻ�^��F|tĥ�h��HY��i���ݶힻ�+���1�YSj���N8 e@t���j6!�̑�e{�`!�Y��������,;ʖ�7�QD� "$�\~�Ȩe�5�O/���#9���^JN*\��"����\#��7��"'�@�0�^7��/!�� �%���7�I�Go�a1u/m?����d� ����ـQ�JãQ�J���7���%����9�?@]���(k��tVCSykh�����:Q��e���LU܆5� f�����ݘ�M����E&h}h�C�&���vp^�o_��L���]�x�g&�@�w��\3�Zr�J�!z
Ak�e���#|'���ݺ5~u�G��w�>=�t�l.I� ��]�+��B�P|*��=C=p�����Z�g;��q	c)	+��6��eŸ^m �xs����k_J=3!ͭ�c*���H_;���C�5�l��$�)�E�fҚP$l�a���}�f����-V�![y|��yGG�XR��x 35��)u����1� ��#��"9�̈o�ⶐ���t2���ƨC�������ǡ<��7/j*:�9��k��g��4�4�)���jE�������Y��v3O�f�9�Q���(��ke���`怘x:5������#�&ŧG��Q�i'l��z�Kv�#؊�`�O��f�0w�i
P�8�y�P���zT�g4u.����Ț��u+֤%T�9H
L��<�����7J�w
i����2G�%�� z�4' �F˾ە��42�2%h� �3�&�j�[p
ݯS7���fN�~�衵n��}�66zF��t��g�Qcw����꟥}�`W�
 �.n��]o�T�j��`G�b��>�H�d�/���Xo�;�I���且�8����̅�u�����X�L�)J7���AƋ�a"���"�&��s!�3��زАS�ִ ��B�G���Y�,�Þ�!ҋv���x<�_�5���י�SO8����,����u���۩�E/�}�d�UPf<<��kf{��%wo��h֢|��z� �&T��'����K�%9���ۿ�Ny��b���9�_�Y�	�c�+�{�BG]�#�0%�MC�w�I"�@��1
�}Y�gz&�g2jQ�h�	�2���_��5�9P^�.��?�j�'W/d����< ��,FX��(�n�	�ʉ����;��`6�S��گ�11��[ۈm���E-	v�6��<A4�Ǉ���%�k-쁝���S�٠?c�;mv6��H�~��B���%O�n�2��0"�'���^�4��G7���J�k�@����fˍ:�������5��=��\�z�l��%����W��
���#�tj��1޹ER�,��E]�'�wIV�y�z��b��YE�By=������z9�����t]�o/���ǡ�߈L*�i�Ϸ�ǘ�ѧ?�8�ܴ�btY��8h`&�)W��8�^��.�5k!d	�ϼ��b4�|�K�b���.M�l��sd�y���q����5��s�y��v{L��~�a���w!o�Vbs'xI�w�V���.����\ ���@��iqrѧR�.���Τ|��o����x���ɚ����,�
4T�ۦ}���Z�
Ro�GCc�ॆ������W��{���j1e�:�HD)>��TA����*I�[O��wVT�V�z�Ol�]8�}.h΋�h7/���F� d׋�i`� ��נ��1>ح\!�ԔbN�S�0Tzj,�Yɛ�лȑ�����"
����5�1IF<����}O�"q����:����ƌ�L5s�������&_���̪��Qp/K +g'9r1F�����۲N�.�Z���WS|����I�n����	��K������PQT�L�{YH]�Z��X鞟�^�-Z���@gY-�0��������H�9|(��YU�p�d(|��$i��wlc���Z�n3�e�0��.5`��>5�|;�&�U@6�%R޹�vV٨�<��2��%�b[ҷ�ݛi�[H=��S�.��}d��X���4*��Z���ཪ��n��*�\⦎��b�_"����b�� ��r�a���wZq��X��JKΑE�9$M\bl�Oom�3�d/M��ځ���?Ay�m�7���7"���$h�;�J�p�[c��&Ԏ��5�qJȗl�#�/w&����۹����U����C�%Zm&��S���ݓD'�m4��3�!=�.VB���9_`O�н�٤?��'�uƱ���G[���F����A�'��Dx�cC�^ƒ�`�L�& �r��9���n/���RA(����1z
T�(49T��ɰ�<�4	w�O����h�|�@�'���\|�jlE���aR4��P�Om� I���|p1i� K��t�Bc����o�Rd�15��k��[K�M�
S��/�Uʩm"��Ⰽa��UE@�x��W����>Ve4t#Tg��݁�!���#�$\���4�%���b`t�����P7���R#dd��N���B�7�m���Ғ�0��+ �F�����~6<���;L
S��ǭ����nc!�NI�V)��ph���G���fw�B��ͥ��>���de!�
��X1�4�]��#�7_�IM�.�ն���X�3%�/h�}�����L��e�M=���7E�7���ږE�ݡ�ˀK���b���v�6Z��6_��!q��%t�`�o�Jc�ʏ��A�����p��g�1��y��^�fJ���A8G�
`8	u�##�䉾����91͚�/�6	H<���6j')�"Di��<򵺏�Q�Ӣ�\���#(� �ߚ:���	���'��
��K�]��^%�9[��V�a�=��ӰwUw>��I����Y�������n�Mfݶ���jG:�)�y"N�=K����k�*2v5�ǫ�I+U���ޓWb�e�����,���a��!��ˇ}��R�.��j��d�D�wP�{�^y�F�7r���������UYѧk'���+oի�M�s{,t>���q���#G�����eH{��N7rA�`l"���|��moi0��k)�N�8�ۀ��z�A3���E�Fdf��Q9��eD��H�]/5H�=��v�f�Lv���1O$�Y��3_M��NbS�G@�c�� �{�.�?�L%Ӝj��w�R�-Ъr^S'\U�ߵ��WH�o/	�d� {�L��
C֣Z�	�E�mQ�W�*�� �Z7o���׮Ī�]�@���W��$z|s_b��wC�;&�=&?>�zωmB���Sߍ�'�s���/�Ƞ��K5C�1"9x/<'�:9Gl!,��H�j	*U]���Tߔ5�u1��h'#ZI���� ��}m0)��e»��'o �r�#�/�:�o"T'�b�'�����VxrT�X��1��<n-��w� �
T0�~��ɟ�(��H_���3���VAM�N���7��B�h�ί�C���C(�?]�H�ն0-�9ۙ葊V.A���ߘ�7�}'�}�a�������ꊏ��l�8AL,���������s8.��5��������~�wQǝN#ÁY7Ae�`�������ҹ�.m�A�`�����Ј�*�m��	f�Ra�w��=�n?�m�̹�iu��u�����<������C=�Aս7�HԵ��P�I��\a ^�_����+��K5�+uEL��+C,� ٙ
�����J����u./��a��[`��Ta�D.+ ���ۮ����U�I����!��܁�J2bЄ�������֘����1>�h9 ���<�\���u��GQen`v��6�T���2f A4<'S-�%kPX�����R븵�E旲�&����K-��\z�7O�8�$%�|V��)Q�P�����߻���/����iZ ����}^4N�"�j����0[av�ZT ���a�K휪?71�rO�����`U�`�i�d��h� �(^�h<�^��$� /��y�o�E/X��45@v�3�sKt���&�p���ԅ_��+nf�ױ�]|��$j O����ݢ�w%���-���������������$0�H�ٮ<T�a����u �/�i��Z~���_؄�(�����,��*1���HEJ_�$�l��~Y�)��==EQ-o�(� 
1�%�O��Ӆ�(��������Gg�1�K:1d��8O����X��4&��c]}`c���E����Uh�8���_p�#�m��W��20h��;�>�ƂS�^-G��[:�3\ ����r3�.})嶀5�tZ��J#�HG��`��V�>졐��1 ���~#(�M�,;������z���a.�ǘ�C��/�n ՝�#Q����@qi�+1���$�iz��7�q�Q�V�Z������\�h�����h�[�F��o����pd� �!d}-tDn�N��l5	~j�Gs,���>V�2��mIc�6_~�fy�7r���/��D���E9�
�p����O��4���E,��H��j�m�?%�e��e�Hn����!�I�'a�@
�Ku=����B#��A��^]kV�������ߴhݎ����n���Q%�ʗ�H��QQ�:��%F�p芋`$W�������Sf1�g���(R1�[�a���� +���9Ǯ�k���ǒ*ɾ�p3A]CN1��|�6���������Ⱥ�6y��"�Z�k�ݝ��A��A,*�T{�Ϙ�9�@�ˉ�5�0wC����eQn�>.w�z`iQo=jg�#hNI�m�Ew�6�t��_�gl-�Np����@��4\�}��8\J�|z2�2������遗�O��Ңw9�aD	Aݣ��,�:G��5ʡ�xID7#O U˳@��7� �4�C�m�P�~j.�K=K�,�{	���_�z]�v�p9º�
�E�f��XjN��7����R�penx9v?��̟p;�a�� ������)ns]�&@�Ol:'�����d �
Fm,����"��F�2��	�!���w̨�@�V �J7PGr	B�b�S�'���UbQ5p۵�[��Z�֔�4�h^g�@��Wl�?�P>�+�0\���,N_���ϸի��M0���>C��HК���'����,�l5TX��3 �P��4X���H"��3���A=��u�}a�\0:�%�b3��EF���'aE̩�Mg��M,贎��m?�,�ӊ�Wq�ʽ
Va`)�����^�: \M�8���=<�k���,�)Q��i�)��P�z��Z�z������F��{xw�{;*�U��:+Eq3\@ySO5������\�O���d&����_��w��n�i�Y8��g7=���0&�q`=h��r�t�pJ[�qo\="�m�gW�Am#}s�V��6^���D��o�i-�	
�e��LH�V����ac
�:�ڂ�*҅]�,���\�\������IΣ?O�ڒ�U���<���0|�e���,@��Y0�����!��C8�[H����i-����6s��������t��&v�!B�l$��]���R��Y���b��R�w!Z�^�h�@/_+�i��������r���Y�|eYP6������z���W݌8���\���p0c<����-ɤ?�&*�L2LS�?�v���'�gD�Ϝ@�p����|��y)�hR��b�c�\>���*ߪ��2�6w���h
��1͖�\���Yg�P"מ�f<v�����T>w��Kц��{�(L����m�ĝ*���9k�N|U�	� �%�e����|��/�O�ĳ�W�@�`=�^�t0,���14}��)��R��q7�b@�w�,���wY<�����B�"�i$$[�&YO�l˟�������ߕl�M#N�v(�Q]�{LX��-�*��9\�%��:�#���Ҋ_nO�Ix��-v��W������EA3m��\M��Gy>b@��>fC�e#��~�%L���f��r��*�7�3^�m�����Q���h����@$� �!B+K��X��#j�)Ț���������$7�E�5M�4��	���΀�LNp+�ah~�kq�8?v�4<�꾶jDif{�+�\
2(�^�g��ɼڶ㙩xNOr;�,2��>O�;�X�g��&�0�0�𸮈�C�@�r9�p�����G'#�����`�<%���#�Zch�@�&1��A�l��Xs�O�ϻ�ф%���͸8�n9-�uRR�����=G�@�`�Zf%�X2�U�ӀDR��%Ǎ7,��`�+,�K����ΰۘP�iH�'�&Ÿ�
���ɦ�A,^��j��I+��+(�>/�*��e����~:F����]����D��l�x����������Ύ�J�/�h�W�a�`!'��[Ѯ�<���]QF��&In5� u�@!��?;��?�J��z��`�TS`�%�:r˹�"qQG3K�m�_{C߶dbI-��0,8���0����Ҕ�4�64}�Qh&�j"WW�(U�`�GR�d��p.by7r�z��
��y'�FH�$2+O�d_⫿vk:sX�Y�F�*ޢv;������y緦�(��D���"�s,ɛ�񀐱�H��̩�o6A����DJKwBƠ���m�2 Bd�ꦯ��zk���y�uFd��p9:h[��a-4N��o�R?.V�e~�U�������3���7[��5�����¼+<8P⣏Uu�lV�P}��
߽�k2���p�`��c��,�n��^V��gm�Կc�?�w�7C�ܭ��AG�}�J�2@�FsfMd�塵	ˤy�>qf���E��5թ��x~�^���Yq�M͎X���<{�m�$�VX~�����Vm�M'B#���=�P�=(��<4�<���/�Ҕw�k�/ΩԨ!�FW6L�4,�
Y��х��v�07�[hxI��@�C�"^:��R�LG�D� �j)���h�'�0n�Ɩ5��>�Oz�o�9��Ƣ캡���y��&�Y��s���~��'�y���8����0���L���4 i���5�����R����r�2�W��z���Z�{˩Q�
r氁�[�k����L�E�@���qjus�\��ͳqdd����ڜ[�k�F�o�t��Q��j�M-}����w��0D���&�*�OU��9����%C
��ޣ#���B0XB��?������D���S��h���jE�q�]RH~�'�	h9z����i��,k<�<�g�P�~��f��v�Ĭ�=o�.�K���m7
��[:[�^�g	7O�5X�v�Ҝ�#I) ��q��J2�h*%|/�~�&��'���e4�������M�9�?����P a�o���0O#O�ݰa��ЮhNdl�R���Ŏ\}�{C� FTŐBR~�xu�W�@}�DUA�zvL��=��cru�!},�;h�<�4�ëE���U�/j��		��;��M�IG���M�\N{Ե.����R���T�m�kԓ6`G��y�z��8��F*ePΝ��Σ��a�$U/o��@�|�Bs�Z?�ZH���<�*�\��-�s�s�L�X(����zY��m���>����Z�L��f��m�mj�~}��>��� ����:&�C�%�T�*�ƃ����.�=A2��lZ�V�%�)!�=�?�g�)�$4�VX�-j<�dQ��B�(H	���Ɍ)Ӌ��t@h`�9��烯̲�|�\����`����=���f��8c8���ac3�� ?��B���ɋ���1�d�(�c)$�V��E��USq�kK�-� 5��aP|�җ[a�ߎ8hl4~b{��l �gW������U>��}x����x��B���4a�/"�k���1?l��
�?c�����\�L������0����nټ���5سF_��4L��%�p����B֛M?͔"���z>�I��J+�v�P��1���&���{��.r\����N�f��t͞2IE�㠭XZ�e�����t:�/�Oow5P��I+Ú�fZ�J4c��Z�v6*����^���@A��*mL-��@� �ed��\VC��T�8J��Խ��,��$��^�6��[�l��iz�-���EQn�"��sK��И��:���("��`���Ő'Xfs���<n�ċ�׾V�I2�<��@�<Q-��VHl�?R|h���c�y���nw����B�覂�2:���9?\�5�K�H���fc��E�y�WVD.x��,�oP�w�U���̘��e���"�
_�[��yk�f}�HoN��uBz�p����X�.4�����S�l�_9�o�mm�<���;Pz�:���,n��Rm4��L
¢�����.���O�T��
.�y߼2��!�řM�U�i�[2W�$	Xg�d�XxCg[y;�b�����XGG�$�B�����ɲ�\����;�,�Ԥ����<	�e��$	o�N*.�+�x>�� 4H��;ۤ̽K���JiV�Q������F�wQ�SdXn��Kl3��ȶ�>BBC�h�_��ޤ#�Qn�לV����\q9 r�떳�a��=k�W�n5l�n����� 5Ĕ�=`�NU�U˶�V'k�r�V~<��"Q�?a�j�'F�Rşg0[
;"ϱ;��r��Zl0Aj��d)e	�n�SD�>��nV6�
R��3�Q�.N��z�=��xT����*��.R����[,[H��#���)���p���V�U�+x���������	y�,�;Ύ��osp�o���@#3/�W�6L[?�'��J#��b��Ⱥ�-�t��X��Y�W=���.�*��Pʓ��Ei����|�:N,`d�w����w��%��o���!��[�q�3g���6�y\�8�ohV�������i���>���joV��`F��nJ�&3����x�;�fGP��ǐ/U{& �����jtf
�Dh^@X����=��s)��W�����(���+��3*0���#`�z��v5��V˿IK.�裇��t����(��$����k�=�xw�P�Ie�-5UR<�J�� ���昍�ԙq,v�i�ۭ�14��A��(�:���}x��z`�A"ǳt��(�OAs�4qԈO[Յa�D%�e(��{�D���P�F@�m��Is�S�n��R�/��imc�qN�T6�B���\�:9��g�;EV��ԂW��=5Ox*qA	q��K�Pѣ!on �ݤk�Ng�WkV�?t`KJ�(U�N���뛿��+U����lf��Q���G�^���Q*�ԧ��-:�z۲�h8����j��m�a���؆�GN�^y���&W��"�Z�}=�F�ْ��9�fZ-"Fa�?�����W6^���<�2zU�Rq3Q�O�b�)��ɂm-]�}��:�`����lVi;���O���d\z1�?�AP	(m�p�rB���)��u;<�b��p|�Y�j��3U����3���[ߍ�G�ꪛJ����~�]���x�7g����3p�o��pa�
��s'ש6B ���z����Z��vl̈�nb�c.OzjH�/��«�>=P<�hi��H�X��6Cx_o��F?����Z13Ү�e�.�ѯ�J�`�`	�]�	{�| ���m�>�z�Xci=&(��ؒAnU��{�6'�e�^����.U���C-��v�{�8G&�&�;�Cݲ8�k�	�����l����O@�F��|ğ�n"��n�j!�Ŷ�m�v7�`=S\iEl~�|2 댺Hbq���z������%	����/�3>�Ci}ע�+7��'�4�3 0E�aD^."��	�6?��Wd�3�s�;�����@�C�M�O��3>ܡ�(���P_v�8��''�m���K�u�䶷������F���U�eTyr�g���$A�y���h�Rw]��r֊��u�{��(��N��B<V�B��$hI�1���h��eJ���R�+�����qV�5��� �E�ҷ/Ş�,o=�/��s|���g ����n�(��VV��y��Qɪ͗Y��tgR}L�_0��NYu�б�T�`�6C@~0�`�%DyAG7��}@�5���`����ڑo�)�b ��C|�����W�U1bH����#��Hĵ�Q����86��B���DLyn�{�SXr_	���"#)z��A#�9����塒�U��2�B�(q�vF���j,M�.�O��w��$+ߴS�c�w��֏{�1��+�O���7:M�B^7Yr�p��ir��ڔXUl!�^p(���v�5��w��Y�R�@��gG� ���رzWRx5&9>�u�&���D��'\jŁ�F��~����{�D]��7�|����$l�E�p��矙���uj�=m�Ru`��suݥLRZ���������<��F.�;����wm�@#�o2�h���ywe_� K�k�� �i�h)�d����d�4�w�K�X��* ��l f���Yt#P?d*P8Ą�(f0����z���� T����śN��IYL���D�ki�����E������I�.���pD'�OĀ����I�~���t`S���{eH�����oG�f��~X���E 1: �$�s��@�Sk�{8�
ȣ,̙�mQr�`��`�d�h�4Cl)���S-���!�o@c?��2ϑP�� T.��?�`�-c?f,�7�k�� ��2z��x��%��M�݀���2�s�������=�Qo����z����ҏ%}Q�@7~Ȱ$%�jĨu|�z�0�Q��oz�A��k��(ڵ�v�h�m=O����R�c=)�z"1�ۅ�+Rh	�Fe�����`U�E+*���b׻��z�z+��c��5X��eLΌW��!7T��e]N������/�+O�wg$�ۍ8��~���6Y�@#�rL�~0��u53���5�*،b�C��G���	�8m��!�{���z�V4zˋ�L;�M�>�9��߿��v"f��&B�}'�IR�4�=1��)�P����Ȍ�1M]Ƭ53��2a͎�ů���~	�����o0�!l���9��F�X�o�m㌑zMM���)����-�����M�x��%a ���&��:9t�i�!�D�^������w5����W�ɀq��az�oS�D�8ɱ�*hq�T�'pk�|dϚ�;�RLz�t����]f&V�i�K�e�!���4�g,��{��o����u(�
 ]r�[+���0y" ʦ�/s$����q�͏�7�,��g��Pў������¬� �\�N)(� ���QX�,����Ma@�t�>H(H�h�Z���l�T|ﺅ�D:f?�ge)J�GA�^H��AVq`1~���b-��jEÆ�ڦ��b�U'�o���������"������N�w~�H��6�r�8����)K�=P֡Z綶?��"�4���g[����y��'_Po)��%7���i�,��3���:b�dʾ� ��,��AK}[K�(VF�2�9�ZXs�
�4�r)�v*��"k\��pc��Bu��Q2X�/B��m�@����@�yN���6�����$��O���@��-6;�����m�ʾ��x�ę�h�y��M1�N��g�.L�c N�*�,��� �1��uP�~�AR)v��3��g]�Yʑ�����ks�X�GR^�+�CQ���$�	V��j����<�_�͜�]�gƗʺ�qW��@Ā��qv�ȷM£B����A��9 �IMm ���LZ&���:���P�)Ź����a^��c�6����P��ËV�N���Ft�x��3�L;�8d�79�B��:���E�[��s��픚X���@>P�����FrH�P�J�o�����΢���kH�?�A����5]$t0֥C.��*��x�Zʩl/ə�K��n���[_�����k������S)��=t�U�o$7�%���yY�J�y1QdW1E�ܼi�t�����8 ����WL�=e�Ӑo�s ��C��GSR��)L�s�w�}�_2�-��������:�����,*�x����(�&�� 9���"��<"���^�?� a���󪺜��D�BQR� �����D퉫�Җ�P��S�۱���~
U~	�w��i�W�4@��"�;|G'#��
bXҏԀ�
�d ��vM��ha3��=%�����q���	�Ғ7䖂���.�Kg��)�0M����2����L�<�Q-�c�5�T����Æ��_:%R���2��"�l�yı{)�;�'���],�9]l�K��{f%`��S�<{�M�[�{t��P�u�l���i^�ׄ������+��|dM�Ӣ��pϘ���a큠mt_ڍ�S��|G�aD1���Z��'yn^\ڕD�dO>��H� j߯�70��H�/�k��eh����5��ڀ�SiS�K�	11*���6KܕQ�����!�'�Iv]ט�b9����J����"�� F|))�~$�,�M�x(w��Ż� ���7Up��H�VMli��"(�kIԖ����r�p>k�LT�EZE�g>NZ]m�
��iw�,lY�Nޤǌm��q��bI���T-ؗ�;߀,����������>�l[�:]&e2�=��P��,�C�.�|�9QَW(� �{~)���\*�����R���(�����b�Z���%�k4�4�勔kb/r s�r(�����8��l��|�4�ԕ+���s�^=���(8]\��ν��Q��[1>HuI�$����� �_7�i��#����i�gtI^�͉Î~�܊�zT#j���f#W({����})}��J��m��I_/ֈa�+��	�l�v?K��[�	����5�6�����{Qh46o�&.�~K����O��ݰ��qN���4\`4�KŶB��e�}$G>�;:nX��XԀeþ �B��z^���;����k���z'/�ssLv�Y��59ف��z����Fm>�f��1�E�c�	^7�'������J��)9��m�p���0: ��zɑS�s/�Z���#�t��3��r��?��iSm8���=X�/���,'N���2��v|^N>�T�|H7�Jfz�(�%T'�ʛȿ�Ŧ�����Pj�/bm#�,=��E�Q-��8����u��;�KP�����S^{���F���������3���ř�h�Yr��\a�8�7�������i�5�_?v��89h(D�%k�-]�	st�=m��=p{,�N0��V�O<S�6s���#5 ��' �FQ�4v������D�����!�E0�\��� ��d-T�p��..qvl�XU���E9ݹ�~��i�e�9�?oH\�ꯧ����f(��q;U�p����ʠ7`t����]�ɴ�乑|����}�@媬�M�X����%Sk~4�܊&1�5�`��2���ލ%��ޫ��e��[��Fhn��đs3Sj]��u�Gl���Tu����p�7D����u��Kk��o�wm�-=X��/�hj�hp/2��.�l~��ڮep��K��;�u�E�e�py���ALB�6��"{hz�a����R&���
�t��̗]jȫ���qxp��=�װ���[;J ��e���F1�A��\!d8��I=n��\j�z�y�S�^2C� �p9#G�0�!]�-Ep��t��1�e��Q�e�8���3q��&@#�L�c#\��
�;�~g���j��"����;NeA�<���"z�x��n'�cOk���Vas��IDƦ��8m��_��g��İ�#,<�����rU��V�~zܽΒH�(ԣ
�U���Y>�KB�����l����m�o��8���NZTX�B�p�mA��BƼ��}ZN����5M~r�N��4�:Ue�`�'=��R�!s��k��ʬ�ʧ"n�mN��
?�iMv���:�A
4QQaFҩA
�B))�'���o��T�V��Z|��`��R�=AJ��2w��E�1ӝ�YF��}�V��*)������f8���9��N�d�@��ޗ�4?�����4��Ů^VОGf~U���n�Q�rNqF�2M��+���H˞$����
��&)Cz5����&�|��:M��Xfd��,Hsy�����t6&��bT��~�A����0c Q�U�sr�]�Y �C�/)��W�ه���.~��	�O��to��t������-���.Ⱥy3�`���R��)3e��/Z]_��cP�7����`��n��z!��X��Nn��F�K?s�@H���/���z��G���dD��x?�G4.�+~��s�	~|��z9�X�B!=ji)n"q�1/|��m�.Sm���@Y�'؎�МBHpT�K�L�-"�ܟ����]
;���'�[�d)��4Rv����e����:m����x����}�&.(0n��/�����&j>� ,�S��`���q����C��vQg�mc���+��������JE:�`���Xvߵ�Ą)['G^hn=*�>IAz�&�R��s���ϸ5� (Қ�qb7^��ئ��Å4��+��>q�}�?q�ݭ��׬1�I�i'(�lb��Q��00 ;=	CΓr��5�S�x]_�4 �'"4!�-���<�����U�ڟ ���l={��&���}�6MT��9�%�^��M��&��o+�����G�����h�ښ��Sx���z���]l�T���ԛ�V��4@L_�f޲'srr�F���VG/C�+i��Fs���1s3TT͝��W����9��C�����D�TtT4w<�%�R.���Ԏ��<� �R5g!�3=���?� �����j$��J%�
����W���z0�D�G��w���IzIM�k���'}m�{�◘ģ�R��b�8=�R��&'4N�Z7�tE66C:�h]�u�K�2w���mw��B�D�%���G'���O��Q�"d���������#�3�RP��!�'ͫ��!�?����S{�ƿz��q�d����ѐ�J�S��g�b`��g�-�����U��'.�[��C�����F���sJjd��&�D����B���1�(,UXܟK^����P.N\�y�өc
۠h��߸�8� ��[OP~�a޺3���p6���1�k���rۧ���߈Ϻl�rhS<X�!;)�|Z N=�N��ҋ �O�b�|���|ZX������+k��ӗ<��?��KL�^�˗q��a2���Ҙ�[!����O�&n��x�����a<�H����fFv` ��� =�Md>�,��@��-�Y�͛wdi޼&ѯ�a�>�������MT��9W f�t:X}1j�`�t����_����C�+�+��$�!s�e��sY�C ��s���ϐ�nd�%#;��u�0�He0�׳�K%Bc����]ĵ��uQ���{)X�{Z����,V �F�������3.՜ɷ�W����;�0�O�/5᷍Q����(j.�qZIy�L3\����Qա���vJ��ӧW*�B-;AU��(9�\r��d�������im���E3��4��Z���d�~A�$a��O;�A8s!���V��ZUD`�ݪ�}�i���7�\<������=f���3X)��7�^��2��~uZw���.�r�<#�K���Y\�0��)cK�G]�A�Hvc��l�*��d��i�0lX/߾?�œ8�b������8�:��ޚm}D�+�^���^ J� ѽ|�F�#^�<D��m��u'��0Y;��&=�m]�!-�)	��ps�����l'!�t��7����UZ8.�Ϡ1�W㖌~u��[�O�����a���/�|G��"%�I�?_)��eè)+@X3<�}n������9���`�q�Ś�g��VKƍ"�.T��P�vUM��(��A�f
�L�������	���̪�&�T�R��Rm�;��.���F��gᡭ���}��&p�jW���#�
�E/R�C�?�E0�W�x�9t�dʾ��}��:%Kd�c�o������o�lK[��ɦ�4�T?��H��bz��]rT�Mu!ք���.��XO�]�����v>l`���eҴ� ���+�
4�G&�D�N ���qzV]��.�¦ ��lq��0W�%��@G�:ib�������f����6�rv�B��_�/� N6=I~A}{���ʤ����p�Gwy�� ��瞙�]�Rb�����͋����K]�g��{�>z��x�O>7���NL�m�'f�, ~r��$*o'�}/�$��S�*'��g���΀�?$�T�#�4__�jȥQA�a2w���ŭ�_�0L�Z�ivUh��d�X��5��BϽ-?8GpB�Ms���C�0[/b���b,5�6���c���zT�?�ȡ�:��;~����{���֬����0�T��}�c'FP�άi^Έpu��ܛ�������c e�;'8\�������O��� �c:܏���7��_���,�*Fc4P黁���� "�,ռ�7ף�!��N~����j ��	��Z-�/���NF���0c-u��SV�l&�����ib�c+o�O���铊P���
�<�W��ڏH�f*���p�Y���y.�����O�Ve�~+L����j�l�Ɠ�e��X���{ϔ��� �2lC�B���B�:
�7���1��i�$���-��T{���B�e�)��py�`^,���܉JL���j�
��m��~u�fod}*Kgq 94�ʇ'q��=2w��=������+��{��KL�IRn7$Hz^�9��V�9j8�<�qQpV)Ps�w�j7(Cb�5%G[�e��R]W�I%��,����.h"��p� �6���:LR���g<C�,��
)�T�|��1U���9�Ŧ$��������t%�bRaz�K��|0�hj
���g�Y@�3�(*>�f���mn�c��ϟ�p�MZJ#������3�
���o�ʀ�Pr=�%���~n��7�j~E�&�{���� �� ����A%��]�U2$�����֡��*�z1�9��C6;ic��?#T�ڻ\äZ��S�'4'�׾��P �nďe���N.�ډT�L�[ׁ�I��?�R�a����z�9�L-8R<B��Jb�㛥p�I<x\/;�����hi"!�[?;�~o"d�֑K|��b��ĸ�5ʒ���Rp�����22#�ysO
Hux���4e��R=P�F��`�]1Sgӻ�B�IC�^"��#M�E@ƍ1�/�M%�-�˸s�I�\�s�N|/���-�"�ڢ�:�����y��t߅���"�Y9e�ﾾQ���s܃��������;Ap�����.�vp�	.cN:<��)e�Pi�^�+�.�����z�fV�l�B'O��Q*��0^��G�ۻ2�~Od�3r2��ĕyRk�Ɣ�\����\M��b�BV�(�@-p�(94���?ğ���qk2S�*��� "���u��*��/�2��}���_�N��(i`�a�a4u�n��w�w�&�����u�������w9:Z�a�8��C����ϘJbԫ3��G��|�hg� �����?��'a��J�F�P��%�yb/N�2�� ��'Ь��rt�X���Jd���o|�6E��׸o E�!1��QXӌ:�9rP��}�b<����
Ҹ� �9hdת�ĐX�V}�A@�ʨ�Qh�y�C�6E+Q]<�-�f$��[2�)wDжi�[�����mtE%s^����O���A��j�m+�U@�m8���l��/4��ł'�o5�l�0Q7�EMp�;�*H�<��9�v7���I�8�ׅ�l )�{��spma�������"ٖ�
]���q�zs>�$�-�e�r�'��1A%]�ؒ��G�l��W���]3�wv�6���gf�&>s�P0+�C��>�7�B�GL��F�,3��ċ���z��NـĞ���;�hDjJ��-pP,L��vT�{j�����!fYB�m�>:-����F�fg��eR6���.c~�*���SwĹ��wF8~�8�?e6�V���-Z�M��Ew��ږ;@��	��DtIX��S ]�V�*P4�1�(:9�яL�����Z� =2����Q�#;0kt���i)��D�sL�\�]�f���	C�ĘA���=4��*��b���o���ُoe]��xtarX� p�G��ON|-��K��29%
���ӈo�Cw}C%�c��
�#0���^���� �F?��\Ml��.eP-�Rw�"��,��><	8\~&��F�dh�����,4FN7/�?�x���ڇY�
G�꫹R�M5v)��n��Y]��#>��W�\v�Us<�^ o���b���m�r�H	e�fj|�/D,\r�A��J�t6�D��������^�~�"��4���E��;��tu�|���%���x�����C�>1��a�q��h�A�ql���+bۀ>�7�׈�`(A�t/st��:s��m��\�[a~�s�m�|.y/�wS���l}ڻU�S4T���;��J���s��p�����W��-�ei�/�Nl�z��oB���a�:�ty�YD��1s�5�����
�����s���A�!�~��������G�������$Gn������R����o�zdO_� M4��3I~c�`�����ơ��S��e���v��<�/�l���i��A��"H��y0�ѳ��0��'���|�-U���n�b�K��O��:�b���\+d��� ���'�A�E?���#�eC����n��� �|lߦ-�N'�Id4<�{]�`���e��J't,Jm�9лc˘�Hm�hg�9#�,A����dr�pi���!����ˇf����W�\�cK/ßb�}��-�;F��䉆(+���������O�e��Q������$;���"��K9�B�2�R +�ü�a/�� ��G��T��9ʪᬫ�s\��ɂsh�ze���]�ӓ�q�&�-"��J)������Q���d�"�� ���?A"�u�{�����*^�:�7[n�u��+��:�U�IM�.��>�%�����7��q�d��6��!o�r>��!H7G����ӡ�>l�.�ա|ũ�#���8q���4����L<*^H'� ��J��5_�z�L���tKQ~Ѷ�˺u����s�VL�o�$e�^����L�qD��@�:�}��E5/���=�:����I��"!9��&y��z�ԕ?���3��Gff�Ȑ�{�Hcfg������V�jQs�2��=o����r�eK��z�wN��'`AΜ�Ai-�wSL�Wz�z)�JD��C�+��C�~�AǼs9���H���G���h���������P�z�ti�z=�����r: Qٸ͘�k��UMGF���ۙ8��66�'`C���~mK�qukia�W�&HƠtSA�ͥ��74�n���{��0X�],��U+�Ŷ�d`�<IH�[y�_$'��lɨkOF��N�f�/��Z�DQ��@�6��.���u�G��z�!�_{�T�����7��O��������.���νa�hѣKwuљ�L���`�WZ�/3����Z0M��eW�^�n'�>3���S\�����դh�O�ѱV+!��g3�����Z��oT�x�Ԗ��-�#�!,���*QM���6��9�:���\�p���o,ӏ�� %o���f��y <QU���1��$W9�,NV�YT��7e�B;��@L��c��Y�yK�N��������/9'�Zi�k(��ZZ	�&.�(�1��W��1�W{c�ܸu	-�_ ��͘`x6r�M�7�n�9f0�a	�Fo)��N2��u���3%�{��GêC�_*<.��j�=W���@i$��+��Km��n�����W�Y����$�(iU�6&o���C�F�E��Am�\�xJ�ko7�mR��/�R������L�g.�t�"�P��,�Y����64�ZV@�8���Z��Q5ذ<����~���/P�(h�/�ȁ�Pb)C��/-ya.y�u~���*\[������.�=	��O>��1H�l�xI���G���JC�i�C����� qŗ���A�!�&�ǲ-+ %?����}�ua>Ԟp�(�-��n}�8H�4GG�5	�Y.��jGC �>J�I%��c}q����Q�[�<�2.XF�`�JYY�\lr{�D:�*72����h�ݛ�g��3q�D��6Κ��VNs�s&���ؒP��'���^�m��`���Z������=X�M�����9H�U}6偓�!��Ȉr���P/GJ �VE�ET��c���P�Q�p��&׎ mR�ϻ���/�M�e�Z�ҷA�|�	C���X�@���o�#���Y5G}��ø�`��-D��f�T�O:g�eMQ�9���3�޹�����|ѳsG�t�(U�I<�QzSͮ�[�n�H�	tK;��d�B��$����)�O �Dn�̓���.�\O� H57���~bF�e$��p���F2۶�3�O�y�J�3�d����#E�Z�K��a��%�[;&ӫim}�*Y�J����7$��AN�3e���N%��&�bE�"����5&�!;�QN�
�}�3�ց�a�E8P���a��"��:c�[L���e̳@��Q$s�^��="�h�z�Hi�)A���$(J;�����g}���[�b�?�6W8�0ӱ���q<�FZ��c�{U.��A���?
3�T|!�ugY��� �[Ћ�K�)q��N$d��ӭv�;D����y��.�������\$���%����]�[Ĩ(�Lu� 8���t�UY�y�lb�x��.�OY\XoX��N��a���Ğ�&*\����Kʳq1��xvE�ki:��Z��G�f��ڼ��3LF�~�n �ڲ�L@�n��1����ت)�U�B�HA�
���w���-����9^�{*���|��W�Q�7�&v3�x�ovk�B5i�7�]��_�XS;��
W�a�ts��ot4��nm�~TD�K��+�*��b1!�O����N���(uR&-�׭��ZҨ=�{_a��H���Q��V�M�0�|r[����B�*��Np��mp�����nNdC�AN��r�LΜz�u_�	�c��KdH��&U~���*3�=ors��;Y�h��3�d��V-�|Ԟ��S6��T#!����Xr��7��kV0.{i�gyܸ_�����N�Јm���	6@��eAqq�z�_�z��Y�>�AO5��+�h7q� Pv*�p�6��J-�
�������yO�ξ���-��cǡ�&�5y�CA�NG ĶqkR3���5�g����P���j`t֬�����g|����O#h������&I�h��?�TBy�?�#�z���	��l�Mҟ��I�0QF_��r%����4�+�����ZC�����Z�_�J���-�6��x�8�3a���y�ْO�W�]��)���5�ç=����/�����z��D7�"2U��j�����5ަp���nIJse��!SqF�����-��Ət3p��z7�MfO	�O�8�ͨҰ���T�Y$$e����rE� qega�$z��BW�4��1�6ↈk8�����	)�$�8ҿ:~�pTͩ�9���*R�M4�[�h�ǆ��:�3g_�}3H����W��W��j�9�'�������" �'��6Ob�"^�u��%"�K��?v���}'۞��Fq�4��%[KG�	� 9\��4��DS��'Pu�I����_~��z��4�-�_�lҬ�I�)��5�5^rR��m����M�4��\�t�R�%�]A��	\0��O؊�~����~@�o��KrSR�eg�.�p/��1��mX͂K ^4�?�G�� !A�y�LX���&�_{D��M�v�����f�0z8 !+>M{V"��$��<EV��Ɯ"0�G�t>8;-
`��;�m�<���\��u&V�r\��ih%�nV�l_�6�%�2*�e��{��g�<���k�[�yY2te@��́���ِLRYd�U�EB� 0�#Kry~��5���Fo�8-��"V�t��P���'�\���U8Q]�0�n�i��p�/�37XS��3Gܟ��� ���IƏ��޾�G��[�!���6w_{�7Ñv�N�0���e�i�$3�Eԅ��3%�9�6߸,,�g^�/����	��1��]�=Ý��>b�M��ڑCN0�9t���f�D�H u_�����R���v����\PY��+OWB{��	�7seԦ��#S �u�)��Y�䕦N�m�KcX;*n-�&k?B�������zg ���i��X#]1d���͇����qh�^d%zt%��<���0r0�Yv�\_�Q���l�Nu��mc�9f�ti��Ke4�a�y���CM�1 tq�5�ޒ�=5��s-.n*������X�|0b��7����b�p��x^��dђB{��?�J�G�C�x~�5r�훟���� ���78T����ذ:��xj��ژB���?<�x���R�a��UbJ2�'�340��
ׂ@��R_<璢����f��!)b�3��[�	Fj	u]��Z��ԫ{�t�~R�\K����i������Ph�b��+���~B�2���* B��$��&��y���P��p�=L�w��s$�ꔸF#؁!O�g����o��uƦ��e@��}�v�w�>H�f�LZ��Ed��yg��ݹ��D�j�7�%k�>jT
߄�T��6'��nS�V�=C>��x����_I4�gd+�e���~����Ok�_X���U�R*�!��e	���cF|��O*U/�kÂL?��xQw���w���� ���Ӱ�4�/\x�Iu�c"g��Z�xa�,�v��wh�g��Z�+�^�2���SQ"`v��"�֭�/�l���N������V�˷=x��*Y� ֗�Fj���݀�1���r�b7^�\ûJ�~�n�����%�nS�j'�f�9����	�y�ߕ����G�������lp�����j\�O��DA��$V�_m��� ���]��76e��;�A�Z5������>O,�L�����L!i|62ʸ�SB�\�*b�Wm�H{�3K�Mt;��/p+09o����]3����L����XB!M��͕��-^y�l�4I���qL�j �A��U<��? �;��N�(��= �[L]�����$���s]�N/cW�?��uh��8�|����%4�7�{w. s���jp�P�+�c�fҸm	�n�c.ZGbʠta���Zw=������;<؛4�1b����"� y�
{�t�+�"<�X��դE_�d�J�\)�_�AS�����c�1|��@j-L{nC6}{��
���t�Eڗ����,��u��7��&���)<���]�V�7B �F�!.EK�R��Τ$O��e�8��C��	�x�֮��:�?���E}I)����8{6�k��GL�
 �2<�sґo��)�nV��Z�D2���1�d����p���E�{�8i��y�#�F��KR(#�|�'j�'�5����IRU�Y�����dr��0J�g�rX�׎���	5�-�%�%�ݶ�0��H�󯶗>T��|9x�ᓇ=����Z���ɣLO�U��z�r��vNw�JiP����}B6,+CFy���VQ�	P�kȗ)ơ��ᡀ�[�FWI+B��k��͂�.&l�hfΤo_���n�����d�㘊��Q�3͚j�*(��� K}��T���ˮ�kN�y'0r��Ƽ��h9Ldt�z��C�`SP�@	b�D��O�!I��f
mV�N�	+w��=��Ą�w�AƋU�`
��(��
e?����WEӝi!�z�z�V�m5�V���|��n�Y>��K�26s]�ѣjv�yide�6MxБw��:��\xt��b���	[�����G��,�-���k�U��e�g�.&�`Fe!v�� �s3��$�/���\|�Vu�u8�h%l[(���zEn��	�����3�I�DY�:t�%�G�Fο�)_�+~r��nG㝤'-�Y��Sk���
�zct�4@OI��9w��;~������E/䯶��^>?EG�(�^��� 5'��Bq��q�	6���?c�f����t����5����C�f`63�>���rQ.�3v����:N9��Bj���F��ǡ���q���{p!�EZ9�Vk����V�٪Lq6��f��p� Zb�LJ~Z4t���e�8�[{3�����C��.:5ٳ���;L�Ly��d�t_5���A��;tP�{#K�Nƿqۻ֐ڿ$t�;Pq���	^��ƽQU�RI�`E�z�q	�	�W!EJ��9��".��]ֵ�ɘ�������`�k�;��5Y�Sі\r�ݣ���vş�M��I�>�d�[>�G�����O�M��)M�V��Y|m{,t;�g"�S��fه��)�Ƨ﨎�<�k��{���{��8��c�I'�"�O�	���8=&~e�ƑH��և�߬IB�Q��F	X�u=���d{/E��w��$NO��^��:�ם,R=Y̽(z�P�"%I�3:�^��yO}��t�#���eݥ��C�-? �[��I�;!I�%��Lc�v��jCϸsG5?m��@�s��E
��� r��C0V\�c-�JU�B�_�K�@���F�@yOv8��p���;�'���_��'���FSz��[�	/l��&1v�7*/?���/�v��K�$}1H���	�>4�d��+e�i��Q<�ш�D�D��H�m��6�J��?�Q:	Ψp��e+εJO ��%]Az�ҽLز��ˆ�M��cۼ�\[����ر$5V(�~�\e�|���l�nO�XF>G����V��Wf�p0��t±I���y��ڝA�w��c.�j���8)���{U�Z66�vw��`�Yk��
��5bU�T55��牆�WG��/~s�P��o� :��:�h���8YU���)G%O�t6�|
F��o�t�l9��(߰8�>'	�����d.K�7��JV����w�)�&�>�:�g��>$��;kdm���/����y-(#}d�\8���@[��_�G���R�V��+F�Tɜ#�U���xT�a3��e��y�2�2��4$A��m���&��!œzo����;��q���F���Ŝw���YYC=��,�C7@��,��ދ���٭W��+U�"�E�B�PW���d@�B<�'d�={bd�-.�4�`-��B����eR-F�8�cľ����a�R ��Dt5��x�jz�B��]�Vd���H]��϶<��b^��h׹�m9`Y����k��`W�I��r���I'}<���l�<�<)x�D�25�ָ��#����8������	�ƌ �
��c���F�(d������Sp´d���������a�^�h ��m��%������e���#7���;���/���{ɯlA�}jB4߲�S����'Scܚ��v���g�U�*x�To�6�".�߽��7#�-QO	9��0j�[�4���%@���9�cZh��`٢�
������)��C�.�������`o����}��{�X]��1�ƚ#}}��߫9�6�e��zA��28��ƽ:�nl,��g�
%���-`�p����:wӾ���cщR�l��V�
R��r����x�U����ʗ���!R���2��6�wq�����܄/�y�)�[h���Y��c���8gS��d�y�"~� ؉����3����=b� ����el7�uTp�~=��Y��E�w#:��v����%ۤ@���˥:`�x��^�4�"2�����^�j�_A\٘�B*4��ݳ��k���¤�.����l��uF_��?�a~>EϪ���3TO'��jH�om��3�Zj�W�)VWA ��"7�E��Eg��u`��"�̀���2&�a�4�m^PRȈ��/h��2J�����o)��=<ӧ�(3&���;j_f7l�����4�W���j^Ps��
�����ĨHL���9�n�y�{����sW�-N��No��/pf�z��)Ait<�@�̵[�ec�Gu�)u��;e,S��ُSP$����q������<��V���J�:}��R�E�'@�_�"�����[W!Xs_�d�J��V������=˞��n���ת�,���.�%,,�w��N�~A����̥�P&Z��{	���v�E\���jC��
fžy�>|�!9�,[�x����j4�+2 ���<+A�$�QڥOĻ~�d��Ӭ�)+E�&��μY�F̭�����6��c谐%1᭬k*3�z�}P��sˠ6�53K�/�:���>.��Fޙ)o���{�(#��a�d��e���/��z��惷�ã!�Q�p�]qK�,���H��N<N��{��6�%xP-���]F��i��җ�"���:�}1�`K��Ǒך�O�u��6��y�|��_[�pV;L�|7��
{ƇI@�I)�K��x=��!��,�@@+����!�l2�R�O��+�ꜵ������$� O�`����0�!��(���,K֊K�  7�5,̡�:q��L*ZA����z���珪{D��AMA:I>\3ٕ��;�R�.�]�h�S�Iqwdo���o鐯�$��,~�1�����"��,���#g�D{��M�?@kx�)._ghS�8=]\�r�W���>��/qC'M�&ج�Tܜ�i~L~s/��򪉨����!��s������ē���ɴ7z��<"��ߗ��,�Ch��xC���X_�||>�abt3�D@�[��xV�FS��K�Y�Z����£��@zi�hO��~�lqs�� 7�F�Jkg`~#,����G��;���3������R$�/�?�Hd��穦p�i��$�IW�9�_j>ϲ
�L0�mFB�ͼ$3��Iw��5m�C>�@t��ك�n�<U�z������Q����G��4BHe#��;Y}*�S���ӎ(��6{XC��P:}bc�!�ـ�Қ8���z��]��=o�kQF/�#U;�}$����f�s��Y$,��Vё��A$�q``S���m��X�U�Nn�b<��S�Ѣ�X�gH��MJ{VFd2bAC��;L���P[�K��q������*#���)�d����e�+���d!*gƧأ�b�`�g?,�#�
��k��� hd��Q�?�x�jk#���رF 53�,�M��u��Œ��:}¯��p�h������'����ht$����T��k^z%)�3~c��L�~}ˮe�`�1G��B1�<A�'�皃�M���%O�5� �/L���g	Ϋ=г�����>�<\۬�"�H����-�;w���y�hzX�����.���_��q�대u'��ws����p��t�Vq�^�����~�+�L��;G�2`O��Hn�k������:�-m�ATah�­�E��9r���I�"�'�Ҍ�V$6*�
� k&\��z�#b�|G�[�����Dw�vAd��k��:=9�9������4� �����T��o�X�O��|ɮsq&U��ӽ��hAž-�:��C֒
�X�?,�i��!�m�m~\��V����K<|G�|��
����cm�SE���[@�u�	m��ay6p�0����F��8��Vy�g1x�����1��ȼ`�T9�����/�Pbt�I��Y��R�����4@��X��T%Q[�!�)�U�|���<7qS :�w�#�(_����@�+пU`����<�L䬥9a��,����B��艹.ۚ�#[š|�ᰚ�3@��Ŧ~y1��u(��z21��ſ9�i1��:�!�&<�:ȶ�Np���'Z����Y������@��
􎌄����_&���� �[��c�`#� TAQW�u�uu^���8�1���I$
]�z�p瘑��� |�����%P����_���,l�	K�ce"�a��BȊ�Z��#|T�i�f�o��Sŧ�?�l��L?����Y%�a�t���5p��e��O_U�Jo2!��oh|�^O�h�S���sA�qZ2I�:!�a��t�'�[8b,�s��K��ƿy�"Z ��zB��୽���F7aE6�6ѻMp����ygg�.�\��@D�a�̳��DֻN�I80v��?"DxVi�����`������-�d��r<$t��2baO�_dG���E���u���ƕ>:�GRȥZk�T+�fvP���X�*|������9���DX���vs�������l�ǓC+��������]��s|l�95�H�	���g�n��$I����P9Z".w��W����Xk���hm�j���YԲB�$ �?ў���{%�&���F���d����Ƿ��ym��s������P�}x#��A�s`��*�-�Y���Т�xd�|���A����~|�lݫ�gέ?�~0�U���h�yN¡;����
S�g�������Ӎ����o}as�v^w�	n}f�9HɜC�L�؜�)"-�៬)�_w[��K��$w<���%� Y��I���� {c����]D�|-g]�x �~5���c*"�qh$���H���%6i��@r��N�s�O�-�N�)�a��<�Ja�󆭧��s�!s�g}�y��CЀ�ie�sAQn�/����8,�Lս�ے��5��qw�Zf��㈟s�Q@`���t�w$��Q��⃀We8nŒ� �&t��8sM��$ϥ��+��~�QE8�oP���������5nu#���7���M!
��� ��0s�
^8�b	�Jj�"2i�f�/7d����\7!֫�E���TۺC�rA�_p*��"S+l��(�TE����'k�^��v|c6]�/f�.�'6x�q�/
2P<�(�>{gmY9PMW��ql�ye<�יV"���\&Ț0hf���m��&d�Z�����[Il�rY�#�sD�)�5�1��ҔȀ���~�$ZW.��+Q�/�tD4$�Q��l���'����7�sH�wa��4������:A����ω�>ix��F��<ػ��81���c�Q�}R��1=����@���d�xժ�^�����\���>*U�GK�>�(Q���Aр��
LYF:S���|at�9���t���r�+��5�H��d�(5Z��A���J�ޮt�Z��ڈ��2%j��^4��5.�Z^}}^@�2���k����4�#�1{S@i�����EsW�I�������96��k�M/H�}�_
.�P	0MCf0�
l��Wk<�?;��.���5׷QJ�*�Fy��ȟ����d�9tY���k��7�z)��H~8�~Eqȶ�o���̃L��:Vϙ�!�w��r:�o����s����"3�^�1��+�?�UY��>a�=���],�<)��r9Q[ryi���=8�E
������[B����7�1��R@��T���5+�Cv��*�^ߩD�z�Юeã�r�Ba�E���Pdao��C���;l#��pm�#�,��ō�KH)���XnR�N���4Z�M�e"h�7������`�CUE��!YL,����I�'�s�M�Ǟ��~t+u����o����~�ƶGymx��ի��z[���\�XG��)*+��+:�^f���;�?�xb���Ԡ�~��IB�Mt3�8����c���<5{Жr���bՕ�E��w�}!�lL��m��>l~�uD9�$a����(�'&�����Y׋\�T�&���gn���p*�L�7�� Ay�]vL�e����k��!�,����,���_��'ܘPD�����lpq5d�E���<v��iO�4;e��x��;��U.b�- a�0� �J^��[��i���H��\M���o�����X������TjP�w�g�{�!�j�rc���"�w�S�Xiz?a��$���x��Oc:��ֽ�*������Cxv+���v�-K�Ţ{�Wݮ�"��ӌIr� /�,��Gl6��mFT�u�v������ړ�KX't,�L���)7�~x�]�E- J��֊���"�����6�Z8�|�2�*��4�2������ْܢ�M���h�4�����ln�x N���=�Ȝ+ ��{��R�$>[O4)A�A�]_��ʪxX_[R�*�-� |�)`�})>�̓r����T�m��a���l�_�Y���2CE�s�׀��V���s#)���l����F1���(��� �i��"���&�d~U�VXz����r�ڄVR���,Q���d�9E$�6^؍5A[��]�i��8��1}�z�;������M׮1�y����&��6Ơ�%	���F�8&�X��u�ǺVo���ףJ�Fo�͠������ԃx��-(P�!J����rLk�qKb�.�%�EK��S� �����{?D�㪒5�,���7����4Q9��KVh�6�Wb<�k��ƈ'|��F����J�&�ے֐]�T��,��ķ���჈ᶟ�{�|���PϪz�y�3�)���)�.�	%ߠx~xTp�s>z
��M��$�v��,�d�n�oȐ�s,���Y<l$�6.���*�gXן�?�++�G����[`��;��-'��R�K[K��b�^�\��k���v&IC�%Q$S5�������%[�\?�v�Y�p�7��ֳ�B�V4�N'R)���ٞ�n"���I�Q�-ѫ�ϋ�9 N�T.A��IX�:k�b��`8����Yl�-<��g�]`��Vp�Q����:\]�2SJ�q�]�<�e�1eXu��i�Fύ��s^zT�
�8�����[�}�B�������x+�/%sH��rIn[��+zF�9�yx�Z���;��ק*�'�б꾂��F�uC��1�賈����GnRǓkP�3��;�r�ګ���$^P�'���'�N��O�}�_ $!OD��N�Į��k��/)��L�1��
,��#`G�P#w\�� ��gugz�>u�v����X?*�$+�8\�2q��Cc9�\���=%�ϣ[�����0�o�U�}���/�eR�,��m7z���.���[��.���A����1���*_�s��"���$�8�%}�Zt����E���%� ��DC�^zڒ�a���X�d�ˢ��$��F�^�\8��f
�k��@��6I&Z�L�������񙀒n:�B��U���r\�~cB�ۀ�<��$���mp\V�q?k�����}��u��h�&�!e͍��/遞�ts�z��/�˽9���`3�㴈���\w��S���P��p�=���3�u�977� ���!���K��yV�kTҹ��e�AF'�#��0�-N;<:u��(0]5c���KX����ʁWd����r~���g�M���g�����F�֝���mN.h�,�΂�?�aPX*�g�j���|��u��n���)=֞45��~��k �k TeH�'�5� �t���ˬ�瞂C�4�3��t�)x�$\F\JA2s��,��V�5�أ���/~j��v��&�,l��i3��+r���5B�O*3�\)_aW�'�{mL�Y�?I�KnVynkl�WA�r,��HZ�lJ8�`Q<#��l��
�]L����f 笐�b�F��:D���4=��LL�.�d�>�%7��/2I�lזۣ}R������B���G/-���|�t��Ez�����p��kDs0���G����E뛻L2�ݱ���L68�X�6�2�w��{��c�����!^l�t�Yǳ��B'P ��I�j��g$�^.5z�D��Y��X$���[�MO���\)S�B��"��"��% �|��·���2� �;�*d�"��ͱ���V�$BP�����1���!L̝/�ia�9t7���D��_��N�6�NytM��<K3ޔx���'>?ʎz��1�WQ�m���e��Z�O�����m��z�p���r:��Z�v��|�
��<��:J�hy��J]xQ>��u��ֶD�.Ҡ	�%n�� "�	l�Α�����!J;�.n?��n�����_X�R�=i@�J�.���ԯ���V87�B�]���q��������p����?W�X8Rx���Jrk 2ۉ��������/0�n�*-����r�_Z��:8� K�·�Ʈ*�+22�>T���"�B�����͓(�+`�����p2H����}~L��A�|���i�����8�d�K�?Q뫏b}I��7�K���]9�&���0�!n7�M$��
a���p�~I��b0`>�&�#�0O�gѪ���
L�`_��N&`ݬ:6���D*�I�uM�l��$o`�+����B�9�T� <���z|$���S�D�H�:/}�K�o��P��j���Fr���,{���=�l�|��
��	8?z���z�#�R�M��y�C��'���Av�%W3��V���7��W�N���N�Ū��l��"�5�2�6MK���j�OZ���ԁ�ݾz��*�ڢ ���&u�CM��.��M��w�g��~�i�u�Oo�v�ܧ%����܁�h��N`�^��+��
�zg�
�P���4�k��5�����.�L( sՋ�!/��av;�}��1�Z�z��i{��"�Ö.�fe���1�m��k��|��[�c�����'�����ge6K1B.������8���}rb�d���g"mb�Q3Pk�(�\���J κ�a�ռ<=d��h?A�9$ي�a�10h���ݜ�(��hs���n1�zU.��OW��j��E���I$]�9C�ޙ�� -�X.r�6��yk�~v�h���~ѡ]���U��Y p����=�d�YS�T��ɅU~~�q×K˼��K�~M�'��w�֓���c䱘*�)��	5&��1 ��d��9��+Z='�iȷ�_u�s"VN���ߧ0Z�/'���A��h�}� ��N	�Q�'��&vF�e��g�7?�7p�Eh�Z�a�R-��A���ἁх�pg��c,j��ݬ����70��>��a)\� y��&�mt;�����D�+��Ͳ&⨌��r�csS� kD-G��3��T��sƴS�*�����[��^Y�B��*�;r�.��;�)D^`��1y(3XΌ{Vַ&��w[_�H^���� ���q��[�3r�7��.L�%#^΢AO�b�������ӫ�]�E�:w�����y>��ہme�s�OT�F*!'5�O���>�4�ǡ�1��=�B�C�[r��
�t�]�,Ԟ��Mo_g��B�+e�XJ��Z%���r�~�9%z�H��o���A�K�EYa`ff��^2E�	�	���Ԣh a��=Pׂ>��Y���U��E��]=��.Sz=��r�k�r][�c��c�]��O(k_�BZ��L����D��h,d�&p>�E�i����	8��R������l$�`M\�����L��Lť�]Ϋ��	�w��"2�B^ �}[�5MO&?�����|�ߤ�5ɩ��](m�q0E��f1��B���UK	���UV��]�Iv~�r�9��k��I$ww�>T]~�x
���g0�Y�l��W�� !����Ң��IH�F �
��n�X��cL2.�V|A�LY��٭����$�� ���8�
��.��y��H�lVRˮ����@,��Udj����ϗ���VJ�bQ�����K �I)Sv��1c�ȷ%�Ub��Eɷj���Y٢�>_�t�P��C���@�=�������`�����s�߶e�xW���%��y�A��̮W��)���[R��$���>Sq�=(��S� �hk����	v�@�E��Ur^��EO��ܺe�p�:Q�E���JkK>���L�'�fJq ��~�MGj�� w"�Ih��֬;_��eY;e*���&kȖl3�����]Pb��%X#�O�StE��M!���+�d��C��`+!o���#m�}�&r�89�p�aiE�`<gR�۪���eD?�<���4X�QNK��Lt��8�z�&��Ok���I �Or:� ^���WkX��-j�;�L�m~�������>L��@n2����^��t�I{�Y�'1줦����P��[���3D��J	�V��
,g�ӭg%�:���O��h�$�Hu)�+�����ֆ�Q���i�f�$�s��T��a�g��
�"fT�8*{��2d�{��k�#���狖=�2d(݄N�nm��]�J�� �m����At�T$r�@6�E�]%BI�̢d�#���X����0R��A�hlڠTN�%6�3�z���QTēÿ���w�1�A\��u�� jퟯC�on�2�c�9���7$iR^�J0����	����Ð� ��l�Rа��* b��N�vX2-4E��Z�,�	)�dk����H�Z]+��eZ�m8��$4 �\�zN%�6���v��C]��0�O@�bF�yIº�>�"EW�=܊Ƌ���8n��R�H�"N�^�'����M�	��]�G�����KKho����i��??sà_c��`�Uw���s�t3R5�Q�)O�*���)��$H	Eϓ���bŻ8�ŗ�v.�P!��5��i~��j�y�]�W≋x��i�b"Ra7�>��P[_K3�����b��T>�[�)e����~AQ�\��e�ہ3UL��Ly�Z!qpk���%��ML<U�GF�W�f��NQ�z�W�I](�}�oT(�r�4���jj��H�9�u���>���ڝ��!����1�D���!p�p�_�N� ���pݯ@3��JS��B\=��*�8γ�� )m9��Y�ː!">s��o��b��Y.�\�J ��1`�̦��C�� XL"V�
=b�Ր��m����ۍ�a};�g!⸦�<.߯��Y��WM�VM�^u�D�fw��D�7~�Ջ��;��:�;�ѫA^^�� LKmV�jO���R0��V���I��z��{��5��X�����p=3�q%��e{v$�T�0��o
u
3:^�O.�'�Mk�@`����
t��n�w�*w�'��B�2��l\_;ނ�������^�"����1ğ�O���?2�M�sV� �U�A��8��P�f�R�J�Ӓ��h��K���%�?LN9+��\�ޮr8��v1Ld��J�*�^M�Nf�s�j�x�!���3���ɭ�J�O�Dou�x���Bd{~���Er{P|��d�K��/s|D^�{�>�t�?���Rp8�ʣ���q/��=ĺ� $n~�Ȋai���S~�v	F��6��"˞��%��T��Tޑ��<�����W�/��!��}���Uu�T&dG�,��ߋy��chs�l���(�
�*C.>��@o����E�/��X���K�b��|F%�o�馑ҿ�*OU�AM&\�����7*�4^���Uc�j�(�b̞����zn$������Hy������='8]}��Z�X��ђ?�����0j��}�%n�k�=b��pÒU�}΅��O�j��|� �p]��������W,,�F���X���\�)�zN����.�ҺoK�Db��jv�<x�p�
�o@���:b��HB����"��]L��`�2q�{�� [^�)%�9Xٛ�����'�1��
���E�7�,��,6��eU�@'$ny]�ޟ~t��?�H��Mm�3X2�*}i1�8�#���	e��;';���T�D}�D���pnՏWi��R\j�B?�W���Z���C��*� �8g/�\��EX�Ϟg1=N7���yT�dN���ŉ�J�5����Ͽ�\�J��p,8����&yM����h�ؔ��ԭ�v�c/��E��+N�rt��^�,���H�Z�K�KQ�g�%��ᐣ����1rn���9��xYAb1�|�yM���!E���Hp��v�N}z��xb@��5R���t����Q���?�&��}�-�H�q)Q�.=F�^�V���N���S�4���J�Rz�5��x�MR�Y���E�
c�ѧLD�@���g��xXI`��qQv��-��z�Q���otq%���R�t��n�l(�muXU�\#D�}���h=�y����q��S������m^��� ���T���^9����b֖Z��	Z�>T 3��qg�hL?������}���{�BA��C��a����֏bY�m���Fã�&�żj��r/���w�@v�r�wQ)�ID��Gu�x�خy�, wF'9O�8vؙ�E�q-��K�U��h��>��x��F�U��p?�xɡ�����m�'���Q~L"�R(��_ R�#��.slϖz���A�z,�+c����:ˬz�7Zwg���nz���K�Ӵ�A68��7)X�1.t����[՗P�c�^�ꛐ�`��;�/��WaW���0r��	~�`��Y�v�N��{Ŝȃ5y�*V��2����O<=��R�>A1�BrP��n8ɴk�g���m<$Lo+�-��-�fo8�⥉�M��8��[��yˡ��'�B�Co��܁m<L���K5�V<�:tsX��Pn�c��K��4% gb��~�I�>/�
�f
n�>�)3���rk�(��Qg'8��|�pߩ:�t������#��8�;��!8��4�N��k���Gҕ]g BL�|�b�ʱ����6h�H]���0�ּY���k�9>�?��k�sv*��liS�>~td�:���`4��ZI�db��+%h�&��À�jk�1I��5�B��;s)�m�.���I� �mN�"<^e�����]���E�� ����_�̴k[��P0ȴ�X�9l�Pi�(ْ])sB�Z�k�S;���0�ol?*A`^
W���T��.��/g��(���'�U��h�P,�;GL��#�8��Z�ۯ���������-}.%����^|5a}>�t�^��f�[Y���&���i���[W��)�F��$=cP���de)|U����
��X��3tvG��(�\>3#^�̃h�����kfKq�x��s> �`�t�W{ޅU8�PF(���@�[61ܴ�-��`�UE�1�QZ:�������u�	fZ�����g�1F�;�Q���1px�=�/��k_+s�Y��.UE|'��H��q����@�31P��:�EQAQ<�����{�s���T@D�eC��sOn�=>��!J E�S�W�8O�`j<F'8qH[uN����D�n�O+s}޿[/W^�"��W�� ��ڍ��{�x��HȊ�pbX&7��$�<�H���Ж�X��7x�� ߵ%��8<�2f��mī3m2-��(�ʶ42F�:u�z��򰍟�i����O?0㤈f��]K랆�~�A;��F��rbG0LRsx������I)���ܚ�'�T�gۧGˮ�5��9���곊����%���Ae.�m&��
�GQ@g���R�h�Ӳ���a�Ub*��8m�*�s��x�S|��Bd���F�/�� I��җ�\d��5��T]�����)Q��K+���HDfw����ECoa���5��K+��dL0ҿ�8�Y�#x
C�\ hg���=�������M���r+�̞�Pa�e[�URH]U�j1�M	�]u�3�3:�0��GQQ�d7@TD���>��i5g��Z�r�)��a\���{^ �����e�T��,�i��d�LJ�������Lj�u+�iW9�!H���R��c��4穭��������.���d
�	{~��N�<��E�Ͻ��&�W�d:����{��܏~y^�&)�Ӽ���s|�0��o�Q�;dŶ��b�6v�a�&���V�a��#,��*�
�$r:�|�G�������%6������_�Id^�ʙ^R������4K;�Ӳf�ޥm���D�������
����D���Рʉ��0r���9Vx5�����R��Kz��BV���C��v�6���9q�� ٨�Fc���.�!F�7+�x�Ac��Ui�r�������r�%������v�i�{�Z��o�bccv��i�G(��/|@�FOA��tͬ��ǩ�EW��ذ�v�&��"�Iգs���V��['4v�T�����J_-��Nz2c:@T ��\K�	�Xqe>PDl��EU�����PQ���3׀������.���%-2gb�弐zȠ�`�;�����A%��m�P���?_�a�kh1�e.[cQ�T,0,I	��3�m�]^�.�T���h��q�V�L��_P'�;��{�P�.��+�O����S�'ӑ�e;�=$V(�E�M3:VF�/�uv�u��o���i�4'	J=`t �;t���Z3�ڛՀ�je�_Q��Z�~�Վ�#R��6p�Zfࢼ�|���Vko$p�o%
|�`�[�0�"���#���.DP�Rp�*��.u��H����T�����l�Lρ�jblw�)WE�����`���+�FY����W��ֶ�w��ȖcJc���o�Ɩ��A��T1��������-�]b����-t��/3 �C�)�c}��?��9�#���J�n�{�\/U�w�4�0W���e�d4�=I���!d�P$��vT�@���Ц?�����2��k�CY-d��<�*,�%'Vl���vXx��v^��]\��Iq�݈$��n������`rYʈ�ư��9��\R䃢``�3R�����f�$_�Q���7���uz��pS�+��>���� Jr*E\	��Az������p�J=��"�4G�y'�#���Cu���S�"��^8[��N��l��ɰ9U�s�Ǭ}ziӽT��k|�����Rc���1��)Z�5�X#鑭{i���#1u��i�鍠�妾�٦1� 7�ί�M���ٜ������Ҋj��0�fh�-o�>��F�'��q`�1;���AEv�@~b.��0�[[��̮���;�Q[t��MHvޫ��v����d(#\��/Q��2�#yIJ�����������mv^����9��X��.4ƒ<�=<��0=f��'��̆~�wֈz,��g%KN\Gi���:����,�!\<N6&Ǆ��Y�a?�� �ſRB�ȇ9���U$�K�cܟU A�%�-��wB����������Bf�����<���;�@�|�#?�%��w#�K�Hm]�Z&�.���={RV���Hd�^W����	�bG����:w�*��Wʯp��p�����>f��k������N+���l�ۭv��&mf��o�8���6<�����t�5"��Hv�`b�[n莝F���"ȗn77]N]u���D��i+��:���V�ߑ�t�^�+.kW[O�i{d�T(���S@�B���Uy�bK8B�=�#����M�D�f���tF�#5�=�9<qJ ��:R���r+���#�re�(���}:�T�t�(��o~��e���|�!H �26��dX��}���L��e:�sZz�L�6k�o�Wsq~[WX��;x-���2�t���$S92�K�-}����$o2��:�j9+ߤ8Ä���zVBŎ�Ǌ��$�a�!��N��`-�g��X�Y��k#M�dV�������kp�i��=:���m�r%1h�F�<~�	�����
!�����PQEz�U�=C�G���,i���3~�S�)!���C��_f������(	Cy٤��ܛ�Sm�7���=�Ҽ�x��n3�:=I7+w�
�@�%S(��5�W�x����0e3�ߨ�^�ϟ��5�ۊ>5XgH���˘�)M������%_";̧����+���O�vLR�҄�*6
�xD�����R���Pr��Y&ѫ�z�y
o��=��+B>*m~e�C�9!u<�0\I�����g٢�(F��Kj�Lnގ�iL�K�$�J�������O.�����7�s�˯� fmW��l�_�{�r�f|���@��;�K">5�}E<2=�K��E�|�{Qdx��}5Z����#�d��L���f�y0w��Z{h��k�W̒ @C����a�~��'h?�SY����rFt\� ����Z���B��hl���VO���f���&[
�!��l��bs�q$����@<E��r�cz���IEdSV�=�C�!M����YX�Y2�ʭ���+T%j'����@���]���.�Ʒ��wYsu���Q���7�g��� �VQ-�T0�jږ-{ϮpLDM"�KL>���c��ܯв,����iκq\i7�rC7n�p�AzAD�4��b��Gu��yc.$�o�eo/�8��$h�������]c�\N-i6$��hl293����:�'�VEr���w@$Yf�&J�yˢ�j�rHD�am��xt�+_�/K�5�#��)��d��5�@�/Iie\tx���P3{��ãM�qg�G�����\�vh`�Dg/,���l݄&6�֞[�}������6�)q@��B>� }� �6'�*xӍ���cb;�co��:�K�9<&/�O�yXf�ܜ���C��y���w�x�(����yf���9=���#f��Y�ƣ-I<�������؅�/��S�r֒�B8yU����U±�J��yv�- ��Zĉ����.�E��d��La̭����|S˷3����;?��l���˱�NG��|։y.�n����Y�v�-�٬?ʥ���¿1�ƚ�:��v]�X���V#��iU���:�XT�n�&A�DCF�i��E8�2jX�]�M�Mn�G� YJ.)�(�K>�<�:�n,d���t\K"��ʶdV�)_��4��P��~��h��������:B?{� 5L�����4�3�n��p��AOG���ٓ�\�U�*L�1��>��}~�+����
�O{�~��jQJz��BsC�D=(�.fc���O���a���&�Fm§�ᥢ1o�Ҙs���q���bc�h(���E���Rh���2?%�/�e��&���R�J��^gsx� ş+}���`Z�6ׅ���6?��'��9��#;2|�G�ƨK�y�
S�����jj2���Ɂ�!�"O�n���v����%���߁�ɏ~JcrJ1�g�}�7��#;_�f��� $k�T7�NL���T�1"y\���tm}hrw�j��x�X 률کswͰD�؅8�lI -��[�ϸ)���$ 7(���W��S�R�����x����l�S�ΉmQ����	[ɶV9�0#���}�3T}�������>�v�6�~/� �G����қ��xyeO̒�����T�7���pj�w�>�Z#�t
�US���>�!�{%�	|�O?��q��ݱ.�E��b9����Gj}K�B�����k'��;��]l�	O���i/󦊃���av�,�w�?��ۮȌX©#TmX\�����2�A��3-���0KO}q��K��=F�'z���W��qC�X]X:�.va��=�������D�Z��`�W��J��3��'����6�5y^>��x�35h�9R@��da�=Lp�1�.��EՓv�b��AtE���������ڇ��-(GzCߠ�QIq
���x��ij�(!62�e����D�n��$ؐ����FȮ����U@��l�����3��v�M�p�����҇��:�`��Vb��J�(O�C7���xz�
��@�T�X���!�U5<��Z���$_�8I�{�Z�GY����p�Kʗ���G@�V��=�0������YN��r*�=�C\�6���p��!=F�����	��v5��S��kU��� {망��Y��H=e��A�Cyiuan��D��''Jxp�z閟�P���g�u΂Ej"�a<P�T��V|�5�����g+��*�FC�%���:h�T5�p�'d����rڗ����X���k4��0JUy�x��'2�+DM�6�#��-�� (�o����Q߯@���_���/iX��w�"y��}�Ag�`q�	tb�o��z �Z��,|�:�WS6��m�Ԋ���Ch&�l��n�`���&�e��|_Ia�=z�:@��
��_ҷC>�Ns|���L,��!�����s4���J-Y�bst���̐e��Ӆ��0�\&�Pp�Q6�;{��2Z�-�gӨ�hX�f��6��=6�h`4��B�%�ނs����=�]Ң�ݣ8�'���C�_�sL�;W6��Ҟ_D2.�&��c�T��R�X��}����(�P*`|#)�X;�%�Z�QQ��Ӻw�@^)��N?t�~& �B���4�WXd9��}{����4�o:����)|�e��{L���Kդszc�������E�Z��$.�vp_�fgY�n�\?@� �T�����2�� =S~�Q�`�HD��G�7ZL���K���ߎ���ؤR��0�|:͚/����I_0�}wsK��4�p���%��V��]s5����?A��
��Ir�Өe+�,��|oEv�����,M��"�\���֍�V.���
ݫ><E"�y������\A��Fz=D�����A8�ϕ:��88P��jD
�Z��*5�!�߯2���4A�Qz�K�'d�mt��8d�y)w���z�ѓ?q����k��R��/h0�9�V��\w��7�e(�����Wj�A	wQ��3ŵ��E1��d5M�A*{�?)6(�>T�g�B��`?���$`?ߎ�	|`
�F�uQ���Ӣ�4jEGf�O�	@�i��!to�)D�8���F]�$�K��q�ly��3>>�Aپ^������j��᧦�8�V��V(6���H����IsK�Qn$Qǉ�c�wpI�
���id4��� -m�%NT��R0��X0t��w�B�`h(`�� ��ʳ���Xy���c�����������v�9-ȿ��)k"�4���k�����߶�>f���-�2~b��Ox�����;Ũ?m>���ї�����W�.��X��P��@�����dR+�,�n�V8ɫ�dPgw�~�z���_|����mEa���Gj�IȀ�DV˰����?v�������$�hDÈ���S��t�y*zE�vCL��-K=UNߓ�%3�5�J��"['ӊͭ�#�Ӫ��5G޶�����JiC��h� �I,�����G�h�T��#��2޶�Ƚ�Hu��y��Ř��$��'Gt�6<�����0��Mn����q�|TרT� �Wh���`Ϲ��ۛJJ���&,���(&�~�&_`�>�s�R����EJC�%���?�]t�EJ�'�;��g3�4��P/�5t�L+��;@=���L6�[��n�T��������#!3����r��`��E��m��(D��^���h��%�U`a���r�DZ�gI~��`#�����5& 5�*y#u�D�!���"�{(!p!����|�%�ʀ˪r:M��R�q2�"ӕ���4��tW��mQpC�$�ڶ��|��D�]��B-��f;�s�௎N�B���E{A�;)��e�ӌ�as���@|k9���L�sz	�9�|~*��5����#=_�lAPJ7"bh�kȒ.E;u$���I�)�Ѽ�bL�.Ԉ�?��T�:1�������@�JwI�z�$tu񎄥{����Fx�G<ã��@~4�=}6��Eg���V�8�t5�`o�l!������w�ɰ�M⵮B��T_"�VVO[�#�ҘnTw�q�}ӿK�:����9�P��?�D��S�4�$d�2�����EmQ,�Żdҿژ;t�)�O�7E�]�p�$�g'��y�mĮq��\ެ\c�c�
�2&x�o��z-�a2c��I�B��ڣ�]�
�Wӣ�:����b�Ǚ����;ǵ6���#����Q�<u����;��3�>�!	��.��GT���oTv�}��#�Ջ���?����%3:���p�Q[���2�bm�]���+���^� O�Z���!.�6S�V � KCYBr�@6b��/���J~���$z���s�1��)c�Syɇ���y2�
�q[�nf�R�Mc��{~��^���[Q�o������937$-���E@�9�֐�{`��M#~��O˅V)���x?�_a�#G����)�4��I�ڽ"��Ԥ	����A��"*9����ǁ�B�QB�9����-��z����ǠM��+h���o�� b�FX��t��z5W��4�x��6๚@8�
���\�,��	[z�*e�F�wߌ�OW��f�;�%dg:L��d���쳎_?sE�n�#_��"KY���c�լ1��Dͺ�^��t�I�`$���L<���/�v0��T[��g��dU�$w��=���d܀�IȖ*�5�����q�!��"�y�q)T&����Dm-��䢍*pV�)S���� hVJ|F��o�@B��ᅜt1M�Q`k~b1C��}�g�!���g��Es��4�@r+����sQ�1/e_�����K�G"�����S�n���0���I�;�?u}ډ�O}�5=ӆt��l�D�To�!+�it�O����A�1�r��7�P(,�גO�N�d�+�H>���#�7hٕ��Zٍ�mq�%�~��2�I	?#�펥ݻs<?��Q#2Vށ����`�n�b	�i�0B�̊@���s�v�߱4�h��#:c�!k��]7�(��?�D�'y*��XI�]��� jP�����D(���f�>e.+Dz�sQs.�(3Bt�
��[s�����t]2Xqwt}J�����$���	S�=��0C���G9�c!*Ҝ!��@o����C�0L�^/�.����Z��?})ƚ�X��{�h�{Q>9kp;S��fg� ӡ�{Ϳ&+��l�k�_B����+$R�(oY�~�z����\0��s�,�b�W��GXPP�Q��&j��O�+� �����@���a������JZ4�<O���>WHY�׉�kN/��QN+uE�Ҳ����R� �
{;�����!�������ʄ)0�'�i�v4�_�t�6�7N�F0��������q�
Q�L��NT�?�F3�����&�㜔7*����%���I����%��K�'�8f����gT�-	�(��櫪ǝv�%���+u�R@�ڥx࠷ɳ{�|O%hV�.qsQ�'`����u�I���b.������Yn��X)�m�R,�rx4���"P�E�7�����<��f�f90�nsޝ��.����?K�2FF�*�8J�����˂͎�S��e����e�s/YlFy�����L��9y|#AI�s*�l#���Y�_�+�ܵmUP�*G�n].��^�s[+-n�3�O�v���A�-bXD��^p'Bۢp���K�_�45(�{>!����*x��I�q�x�[3j��<'g��e��"Ag���n���&w5Y^�)�On7��mE��w�X��>�HPဖa�vGa�z��;��,�3�Rrp���(褕�$���O�����|�Z4r׸�.�P�*y&�Y}��8	reL�V``5Fߝ��Nd}�^OF.q9X(���y�	Y$r��dY���ę����%��������j~~g'GX4��ea��IUZ��ܣܣf�f�J=z�!��qGm�l#��z�-]$Ez����i��{��eO,���5�`���l�`�*^m������0H���o�e@n�]�#I�`K��5��%�`WsF��'��Q��i���p{en,i!%���[��xsL�d	��.��h�����$Hz�@x��&�%���n-�����>q��s�Uti�Ql{�����3o�W�;��U(�Z�f�D�>��r�����K��o���8���gF�1��gqh�Y����S竐�Z���K�SC![m�mO !"�Ҙ��[���W%�C6���`&Ja<�fk2��R�ڤ�N��4&|�@��4�{��Q����Q���0�7�KwH��Ou�g^��i�cI�l�]%��މ�ň�k��
�0+%�-S�@�8�77
ȧ'�8�<�EN���&�8�՞���@3��uO�ukZ�\"�̪9��E�����0�.�x�g�LH��b��2G����P��@?���L'��V,��9
(�o�v��B��y4-}n��r���β��kw��(���W0nd����w ~8 ~K}�w�/!��ޥuX+<Vv��*L�!Q/��+����*��Y'�7��0(����	*U�FFg�M�����)s���(V�JF����:۬���(��1QC�c50wF�_�n;�m�g4e~��g0��LS����4�t��qڒ���ՙ�}���}�%j�t<��j��2�:-���Im<�wz[2H���Y�p�d�tB�\!�EN�6���XGt��OE�g�yR;9=�k��6�%��Bǻ�)o)jɶT]Kݷu>�l�*���qn=LnI�@�&k��V(����%�̑��'�Ν2�A5S0Q3��bA&*�i�=F��P�E�#m�<����qzpt�Q�LO�N���D���C���nu�k�k}A�0��Z�fѸH�LE����A>�s�t�|ܸ�v�I��'�29�G���h6���S
���8?UF7���H�&�UH[�̩�F�����I� ;�Q�djS;�"L���W"�������_�zq6C�����95���������1�k}_������Qx&��]�.>���1l��a~�V��s&ş�[-:Gm�$+HO��������A�.�r����^���/��(�(�$�̓���dc��Էdo-V��������a�0?�����CZ)�]x�K;_�=�xle�L����P��qTj�h
��(x�	���^wfo>�͍���7�A֖K�+Җ�Gr#u$�
b�)mF�f�o��@��UG����]���R� na]��[MK�0A�7	3�=�`�����؄)�h
��AJ��q�#d�nD&8+���w4s�O+Ǚ���İΠ�{jU�D�ʁ��r�@ciG[]5�΢�_��BzE�G��G�� �=��'�����!k�����Ʋ��A�([t�@�.��ܨ��ć�by�ȍ��΄��-=W�ftq�n\욡;����qY������%�`���R��e�׆r��	~W��+kR�]Oa*NF�Լ���&_�k�کƚ��4d��$j0���R�5����[c��	r��N���"#����KO��3���1�
et��su���6,!�ƶ7$a*�
y�?��Z�F,���7Rii���1=e���{Q72�9��d�Y�:5ô�w9�N�Z�-r��O���0�t{�g�(�u~y0p���D���B�H�S˥@k�\�h��201�n{�A��ɣ�	3k�[}��M��&�����0}8P�c!����z���42��X П���
�a�Ǯ��!���"��bCr)4nyF0Q�e�L�_�CUhZI�&�,Fԥ������`���Aׯ�]H����G�H�%MQ���}�_����b����7쾉��e�*K�7;޲�A�l����u�H���YO����{���f7�O⊱���ڮ=Rpf~g����܋m��ޱ�䟔�1�`)LVe�q�.����(��GP��FO�n�A6��RA�����y��c��RC��d`쪱f6	E<�<��)p,��m��G�M�D�[��kc��1ID�쫼U�.�E�7��p���	V��o�g�C�x4i�_s���FJh�:M����4%싱*���ob��<�u=��;��uz�	[�D��}�X��K��Ɂ���d2ûF������"�G����4"`H�)�k�P���7C����,c����rn�����q��o�28@b��%r=%��<f!��g�u8�ĤO#g�hri2̰���&k7�Y�u���{ҹ������~�OG��q��7D�Te�|���q��v�fl��Ohz�v�(���<ц�X�,H��������9�r�p̩:AZb@y��=��T�@�+m�вς��${7wܰ��\���d��� ��V�z�@P�N�s���Dd^��,�u������w���P65��ݢ��(�eR�O|*+�a\ܔ0�����y���3�-肇j��A��W���C
6�J�L�r��hn�G6�K�A�Q6��x�1�n�A�:ZL��OQm̦�]R�H��"f��I�J�0i`�*G�	6��c��آa�>|X�wӷ�f+�b�!�rM`#̱g t��로� X���#� ..(�
���?�-_�D3d���z�Bt�OE���t�����x�r�QP]x�+>���l�7F.��%�a1닚����l���vZBO�+6wR:<f��BT����$ߝ,����5� ��x� �T(�͝v��i�?�*���®�i ���j{������0�astK�,uؤ�|�5dxO�@EQ(#6��c� '��:��W��V��"���A;A�v��*"�:���Lr�E�����hyP����F����;���ͽ�S?���
�����׏�=¹����D>�n���hS�	�WXn��d@��Ew��}��4��%�H0�%�H%��#�G���rmĀ
L�A �R���]����YʍZ0u�d�>~O�cw�19q��M;�}��X�i:���qu{�!���j�'Q� �X�D�v!0����5m�C<�$pj�p�O��'_O� �
�a*�m&����'/�(3i*&�Q5 I�	 >��&���Ƌf;��)Ć;?��^���z�n���қ��G�y9"�7_�(Ǿ����.Sj���]T��5�1��A��2�6�p��F8�D�n)�U�R����D��:�gt���nlj��� *����`�O�8����S���^��i\����v���
#V�ZY�u2�:&�!B��+Z����g�We��`�e��8���h��znZ�P
��vVQn�%v�͔��`���V��4n��D�����> s���"C�L*,g �E���3��1Cݜ:�ʑ�\����Q�)Y�m �Wݩ8�b^���i����N�V]k��F�gw��:��"��&�4�;J�*��S��m��G�g'��yk�9�`0�>O@�B��1�+�J��Ѕ��V|�`E��=6�wb�T������54�m�4� 5�M��m�̸�����R�~R��"IR�U��ɡ���4w�N���( �����J+�Y8���(6B?���tn3�%(V�7TI�7��ߡQ!!,Mna��$�b^Y�A�$���Oi��KD�L@�7ux�u|��"��0�О̪cP��-�߲C�0���@�:F8F^��Є�s>�b���I+x��\Eq���[���W<�9��n]��
������g�c�4�����`��J��ݬ�B��Zw��9f&m��?�8��h���|}0"p�0/�wg����N�c`��m~�(�Q��w�溙T'#[�|�@�شV8\n�C�ny�˥�up��+ݹ�gk�5z������'?Ԅ�.�[(@�Y߃��!/ܢ�撼��w�ٿnE�O��^[��NO{�(9�|+�VݢL�w�_[������d��W�IH�T��W!�gN�?���H�����?
"֥.�=�ND�Y�z�����f�\�n#�X��5	�V�[�B}���?ǫ��[_��w�*x�_Ta��)(�}}�
(;ƻ~���9�EU~h�-����SM�,/��b�ۋu�Jo�pp}{:�`�ࠆ��a3 X�`�)⦌�'n�)�a�h��V��g�D���p�iM#l�d��KX�(��gt�L��4�Ӧ�����b^�2#�9uF��r�N�[�+���A.�NFL᷽._��l�g�@.�-8�s�*�P�1�'�ݷz#�?��P��vD���s��&�V��]���k��s��2�F0Źx�8��j֨QG��Q�WO<)�Ш2�]��*�-��^��p��F]��6�?_��0z�$��x(	q�0O�~�e���R�&\Ik>��耏���)�B��[y�$Yʡq���{�]�a�� � e��ӝ��s�ݵ�C�\�T_��P�\���קc�H���V�^I�������F���'���	U�d�Dx�#h�D����o���[���� ���H���������R����OYߴ`7�JV��A��4�dX��I*`X�`�/��*���g��B��������4ve���./�Vg��ڐM����;ZV�gؗ��J{�����d��.��I���y��@��S�R�����ѡm�w�|�k�����/��s�u&���*�ڂ�����9��^�T�߼2��pZ�Ȏ#����< �'2@yM��&���TwƔ�;}�[&��zOs����b��v�d��S�v����hTљ�����s�z>�J����}�)*��%߸ɕ�}k��w9����\��石�G��H�-�5\c�w	�s;6L�'��@p�.�3hE9�	yRd��x�*���FV0�j����&�`�J����
���C�Dg�N��fF?���r�	/�����,y钺T$3S��g��b!�'{�q���ys�7�����Ńxtҙ:�u��Cׯ��W����ױ胮K(������LF9Z��oQ�2bu5;.�$���O�*���D�L��F��Y��yd�)��1�d#�%�է��t(7�*��.V �m��d���~Sqd{��2�g>��'��M0�2ӡ96���*��2D4�u8���;��1Py��x��ݮc�u�����zm�Ha������a�_ʎZ�:�7n��ٕ�<25h���"�Z���E����@$�N��25Sf�t}��I�c4��I[�*{�A���)5oBTM:�I_�!⤍��o���Ǚ��ΰ�6nSXc��y���v��j>/q�Y�����ھ�"��ys��t�P��K/�!~�Wp��PI�4���[���:�$����|�+.��v[�5��-`t'4��ga}���#�zb[���]�ّ4c؊��r���M7����&yƋ��[s�|�G���H_�T�$ �+��
�P؜Ԗ�0�-��l�@�� �r�8����(TA��@~�0��w"��c�H���/�FK����IO�m����/b�E���SaG��l������G}�&7ň]�y� g�"x�<o�*���������?�z]JЉ��k4��LsC���O�i kZ<�\�һq�a�i�����Y�J�
�Uatﴹ��j0�w�zN�ZA�:���E�����ͳ�!,j��O�F���-��=}s����m:�l��o+��J����[�x(��tͰ�5�A�zJ�C�(���(3p	^*JI"0m�e��� �5h#���u�8Hf!Б�����w�7.y���:|`�+v��d�v]%~J'��%<$��g�3�e������#?
��X�V4�4"��1���O+�Z���fV���Wk���9$�2�bs(>�Fï�HE������t�t��Yĉ��i���F��� �Հ�9�����@���}/ћV	�Br�Yۊ$�;s	���޻��C@b�["�NT�����Bd� �c:	����,��Ր�(|�({V��=�2�ş�����k�-�/����,H�i���z�����h(C�m�\���y|�6��������������&2���=��1��y�[�κ�E����
_�>���`�ѠΜr����[�;A����Q�d��Ӎ7�ƕnjo\�tƙ��!9�1)����O+��
�Ba"	��Bɉ�c���0g>F���JZ�,I6ֵ�zP��U?֩!^��@�W ,F.�u.ٵ�Ae�N���
 �-�o����>�-��y�����ior;�p�
���ɨ�j�>�Ѐ.k���8��|ef~�_c;�dk��~�c.݀�Ǒ�r��P�W�=#NX/��q�����Y"�iwFv���0���L|h �ٟ������z��
4��Q�t�7)����\F���'��گT�1�<Ӳ�z@=_��D,sq?���
��e݂��%���O� �P�<Ἲ�%�=�X�8�{�8�l_g䣻xA,�c�o��1��V!U�L�0JhjɜV@�f�4�X������o��_'�;ŝ>~C�����s����w F�NAnp��������U���wx'�r9]9$Jv\����)H-��.B��3����wt���E0�:����.1��i�iB�ᱣ��ؔU�����?�lؚjT�R��-	��=��gYB�3��ʟs���O����(���û��ʡ4������H;��]9�G���Q$�����1~Y��|[����%@���Q1��F�B�D�al	i�MZ�{���&���Z�]v�=ښ�i�'Y���*�@�Fi�:2�6���!)��|�ni�g3�>R��]�%�d�}�e�����WA�Ką�������ؒ�޻I���rPoȪ�7��Q�N�T���uw|PJ=�N�Q�:�pD2
�~i���[Θ͒�Z�Ʃ��05.h��flS@�����(��M�4Yv�ߎa��Ӷ/ۗ�L�,��� �
�K���/���2k;Y�I'��l0��n2��d�2L�E�ׇ�l�4�(؝_hl����y�q��=í�/���k0���MJpC�D��Z9�����e�*pc_�W����OH٧}w_P[�4q����p�����s��VA����3�z�ԧ �3Cv��&����p6:��2�疃p���hmjrf�X�Y*�<��Ŷ��ؤ��jR�ʅcW�u�\ch ��$�*�'��77��1��q�&H7����\��0�%��jy���$�_Ā~WV2�[��[�wO�L�ȧ�5j�f2��B�t&�����flơ���2�}?�a��8 �*�qPi����_o�g�Ě�M0�q+H�	������>��׆��f��9�}���v��[�.;�l�{h$?n��/�p�Пx<��4�iI�<Doy��������8�s����tJ���3"Ջ�$��	��b����:�� ��\J"�r�d�ډ��p�#j����9�)�Y�J��H�����k���{JZ��laYݯ~E�l|z�/�#=���`G���0��j�nv�t����Hj�*��]	���Mx���H�����Ă�cY<�	���jQu��-��DT�g�d�Xa��1����P!'"ZZL�g����G�1�<��	�2��Wl�NB�2��y�������D�4�H�G�أ��&��iLq�j��u)�&�=QM�At�n�yn}CLtg��[��$]i���Z�a���R95�{!~��|I�Wx��.e��f3��%��k���5�y@�ns�_�YNfsC�Z�qcG��f��{��hD��(����S��	��"�x��@���#�G��<;]���|v��(�~��P��k��$�ArIs7���%Ez�\#
���Xx#��|#�O=���;���ĉ����ǝ�t�gp�<�W��[��(��bg�
,X���z5v�sp��2c��v��g4~�Dk�����A�w�킶��E)7���z?����sC��ُ0X���R	aεt�$,���xj\���3qӊu"��[.�SS��tWN�T���LJ�7]p}��6�ngp �l=��.0�3%'�2d~Է����am�I@;'#�x\@вk��E�%�Ifd9�/�pL� �)���C-�}���Ċ�C�Nu��:�K�K�|V���ha�u6�?��,�G���������o� �Q�s��&�Pi�kC����ok��@�V�Z֩�o����񰰼��U��kT���-L��tP���Z��42������	�>�>��s��{U/h��r�E����#?و#����j�z[x��i��c���C.
.:�o�F�P�?�N��'A"YK���VxҜ�yq[ZK�����v�7D�&,Ț�'���c*%��3I�fPӀ���Q�}�@\��Ws>;kïQ���}�`T��V�n�7��.�u��.�'(2�aT���ʌKW�<M^�ٚ�?4%U.T��.3����7ܮ8��	�;V�+�`> {%��6�5+��=Cu��	�4C�����Fy�*�k8�(�AOF/�x���N���檽�Ze!�&�_A���k]nb�ޅ��@͓�^�O�E=��=��kW�x�=�,^Ñm������ძO�ᵤ|��V��� j�m�~�UNi!��!f�×��Um���MĢ��D��F9�0�R������Z�(~��0y|�`�ń���M�)Q%�ǉ"`�0CCQ-�(~
��O9.��1�>�|\%,@����d�5wB��7����(į�<�� �����,��*�vF>D[��P���`�?�zg��y���C�wKc�Tt<v)���M%�R��qb�U�T�0Q�{bd���u��#�,�$�x3Ɗ����i�u����:k�]�n���w��!�V7Ĝ\|�`l�p[��V���Fs��Z�D�PD��'`3�4��p�5��r����ͪhg/��^S�{�K�O?
�I��Im�8�"��|/0�B=���[��SǇ��p���LA�兙C�
#�xP9� �]8�"S6)u7P�F�X�����W�3O�t{�Z|o�#�(�����ҧ�/:*�0��2#8�\ܵjNQ����R�ib+G�嶘��Q ���>;��A��l�Z�<䂈�b�ċ]� ��h�T��$����e��� k��z������+p�U�Ϫ�X��h8�v�j��K.��׈���:��΃3��}�����K�0н%�s�Jw�l�!���čn��P��'z��Yxt�o!���:Kk���:���d�naJ�����@���]���Ќ�SVN�����k�T�357om�=�XCJǡ�\�IN�|���PXs�!izĿ�=O�2����z��t���/��g�_=A�h=����T~�ٳ
��	f�`��@��m�.*��Z�W��(�wp�b��sM�v�C�����\����ms�l�8�W�!'�1/�����O�#à�����)��\�+�� ��I�Bj�,�uL�V���!h{J7��e��t���e�AM��[�K�͏���V40�g��$��5]���G>��C\M�l�R�/����:4BV�8���G�-6�a
ϫd��P&�������r�)ޔ�o�|+Fk�1
GبL9o�!x#W�)^LI~p%IW�ߘ9,����˭����-��~����ȟ���m��ս��Pm�h��J��4�좁�T��,�Py�P��B���cIo�&,萦�i��e ����X���!FNP�2^ONC���o!h�<�ġ��TgOw�8H�u-�,��*��$�/
���q��77�@�N?M_텃 t�n,�������t�:�����Z�t�e���"���@��u�~���������o$JӚV�8;��3 ������8�[����j��탶ʜ�o��(�*��
Sկt�<�E��U������;�>M��&��N[�M@A1D��K�*}��+��H�N��	�ޯ�Y��D�W<�Q���׍�	" f����_ sE�	݀x�R�K��K�t�`𿀈;;CE�_7W����L�C�z�ڟ�f�ƆU8���?a���nM�{�|����ڤ����7�Sx� ���˾��6� h t�>�W�fN��hό�6JneM�և�i���1��	���؈�1�Sh�+������@����D9�[��'�d'��r�͗+���E3�#��l���x3k�)���-�Z�i��w�v����E��7�Oz�we�]H��)��� �`䉯3�R+~�TmE%��2�;:����,�G䍿uSA���Y�h��fo���x�rȸ��f"}0��)����������0�T�u�eF���Tce��ر'�o���h1��-��}3��/_���:��
+ּ�\�Қ�E|�S%}	D�D	~@��n���n�Q`=}7�3�vґ��ә��q��P#8��D�'�b�4�E��<pؠ�!k^tN�cFb�mn���!0o36�E�	c#�:x�øS�))S#�7apPy��z1����.+�<��&���3K<���$�l���l�c�յ�B�Q�4.�e�	�[|���_�#�����JT��ri�jx�;v�_9�`a��3���ߪE	"��� ����'8���?N<���r�)E�0���ה|�YSwa]��x�Z����w3��E� �o���8�
����-eB�t����}%�LXX��0�!�֝ ��^#)DC�eI=*Һ�j-��
PY�MH��*���̄��:�6ԩ)ԻR�P�3�� a�X�ӣ�/�]z�o(��q���5?�ka�43�-��q^ZyfF������*6�Z��.���%X
��^�_�K!��wl��4<x\e@M�~9��6苀�{�&hfV�)�/����eu�� �|U��۠���O	6�u�����*ŝ�sq����pQ�Vv����j�(�hЊ������*���MAvW�3��{�q=�'����M�!B8'����_�,;k8��7�N���q�v�G("+�Zx�ka�1/WZ9���?�,�/����T�{�25�A��J��t$�wP����.�֡D���)�v �h�ul��Z��i�-+g,÷R
ڭprL��@���  =4"e�*i)1���ۏ��R�x��5ZB7�|��S��|�?��h��ͽ<�q��:���n��q�ﮆ�g�K �s�� v�H����ь~�1��Bx�v�E�:�z��k2�k?���ȴ�$W|b#��T��9�������В,�˼�C��:he���s���ƺ'�f}�7+m�5��M�\�u�G��4���=)�-?>���z��Q�A�<���-����l�GB�W��r�񾭛�Y��2��(k]0��ö�kP�7���H�	Ϥ�ڕU��[S�@�՜���O��`�L�V���
Ni�;0�8����ѽ���Ýw1*��juƉR�+��L�D����&C�ⴼ�6W�a?��R���@���y��&�s��@S��؇�T���\��/�"���$4����-n7;�w�.9jÂ�b�H�e�G諜?�s�.zu���:8�"#{0:���<�&BkY�ኙJ�I�Wڿ(D9/ +�o�=	u�dVw���X��T�2S���>�a�<�}w{Z������7�P�H�ݳe羇~�2���X��JO�{?8m3������5����T�`�ȳ��1���5]+*��?�������͐�9Vd?��Z��`�٨��p@[�h[W�q����ڵ����k��E��ώ�y�LL k��G�n���b���h�7��.ε>�<��鄯��и��rD0u�?������s���%L��{�P	�Ƶ�EߞD=^�'�,Z��Lj�of���(�v-�V/�\��H��g��a��z��(�����mk��h� m3���̶�o b%��w����~�%��_��0�`�9Dn_�/a�(5�\B:�/8C��6��BU8x�4$��l�|E&�j�^��5��|ˠ6����T]2xV�K�����+-���ѻ�b-e~��	�&9z0��g:�W����=hE�l \zh�d���i�>�`Qa��2�#\�:p���J�{�F"��,I��6�:�+L���<�|<����|�����8��.�-"�!�S���<��'Q����֬�	��,T���8{߄-9�o�N@��sl�{N�}�`J)HT���٭F�"��"?�ļ�օ�.HN�F���T��IS܀�_������o��q��7)H��"��L�#Z�w�!�����P "�b�����Ж��5@�ӯ�kC
����b�n^�vw���� ����zd���_n<�r`l�x�s�i`�d8���
�F�G厪�%cTZ.���y.;D� t�&.�����;�h�sz�klq/�Qw��R/v�ɽ؉��7K�x��<��M}�����'�j�$z�5�|�����T�|z�� �p}n�J<�Н"4<�H��H�X�R��Y��
����SSM���1ep��X$e8��m����;u@���!ǃ1�F��6Ä\7FY��<ȊaÝ9�����m@�T��v%����m�����y0�&-i�'��ܩaTl���Z���0� )f4h�j��}��X�N~=��IU�۪����w8����z��V�
��@��)h�M�[1���!*K�8GuP]���ˢ�NvP�����0mB���}��G�Tߥ�`���K�<2�a�B�.����4,9�{�ồ��P*>g��A]���V>��B�Ua@M؊�gO>�U�R�9���8�,��	���}��%��(e=Ő$�P#�jy�Q����χ�
;�l��!z@�?q2��f�pU����Ԉ)���޻��g���v���by`I���v�y��f�gW��d2UL��{pc�+⹹D���V�;n�]��uڜ�8�)�ZUf���N[��S<������ �?�E�H�5�����=a���b�"�m��v�
�wvJ����i+L%j�wK��ڝaˎ՞+��g���e
�@F��H�o�<��c��(r[�V�k=�ᔄ��� �Wݺ9���7/�_%���\���L��T(�#�:��4��X@���$
f��'�b��*cCZ3q�ކL����a�D6s7�Ò/��-������S�[E&6��]�,m�����b�¾���f�6Ē.�^��M�)T�*�a&G�K�lH��⦫���Q�f%�N�v��pr���z��V��n�v���=��?}'k굹��T��.�HjFM�&jt�M��t�i�[J��2�X�Ta|Mi�z���s�WA]�=�c���">�ߔ�֑��E5k�����d��2b�>�D��q�X�:�D��b%���,�,y���_(ƓV0ˈ_l��ʾ�;	z)
�*9~?���uo���&z-JmAb�N��򐕆${բ�E�q�R�H��:TdX}�Ҡ1-�Jne��:"B��mN�iU6����7��+ϊ�!	�؅�\�]����j�,Ԏ�q�	�� �<���ʬ w�P8�ig���D��nz��@�6_��*����f����C�K�8���5��O�E%�$�BS+zP����`��0��&��{"f�_�Ǹm/�R�c�*z�VK�4�ٺ�&�՜4��B��{'�/�N(�詽�Y�}P������p<%�˱[�&�$���
���%�=��*%`d1l���4�Y+�U/�oA���׆jX�����ʖ$Fj�l`H�6��`����8���v�E�)Xj�<�/���P���U�GЫ�������4�z#uYr����|��"��%rkс3^��Z�
�?����JKoYOTD3�k0 �_�CF�Ԃ����ٳv�w�6,*��P�H:eA���8�Z��054\u�
%��٩4�S�������(E��}xp�6]�����8�o<C���Y��Ty�K���o�.��B����VO8]�L�.�N�C��5�֥Yk�v"�˥����K?�? :��SG��=���O%b��_���D����^)��I�{�/�j���Hh<�!��c����F�7��[M��\/s���n�ʤ���ύ�Q ݰr���g����%'1�۪���ܢ[��tBϼ��|+�ɪI�ԨQ�Sh�Z8 7��d��磢��ibz)\���b���oA�Cs_��W�Y-��F����	b����U�7�f�\����GJ5���F�K|*��qʝ�b7:���c�qB��fLx�C]�/��9#5-��_L/�O�P��?�n��<Js&D�4�묘�*��� B0�r�vh�'b8����z}��@�xKXO�\�#�9B={���j�(�@ꌃ�P&��"����搵A{���RX�p}��?��8z(	R&�Bi$��(�>~p�����G�Tib��ɋ��`2�gc�S>�Y��'��u�^韜����V|N��.]"��}��s1�n��C@�S�GPz� |9�mN���3�b1�\!�iqR}訓������˂�/��u�'1XXk��^��"�v���:'Ć�5��IY-r�O�ҹ��K��{��%~+�ff��f���+ÓJ�~��H@ή����Pb�*m�1��oiȑ�����tI;��C��E� u�q�92��y���v��[ ��#s@[��Ӥ����:0�[��4gP�y�.;5����3�����6�'�O7�|�����jF黴�n{?~��� �\^c�,d� ��A�+��P�D��h�R~O��g�Bg-pPd�v�9�R�@Nȶi�u��x4�r�aΚ���-��k����kg�"�K��;�~��G&E�ϠpZ��F���\qr�P��s�F����M���˝��~X�@]��V��E�:;-�X{0Eܾt6�Ã.nu���_(L��[����յ�5��Δ Գ�H��@<�oJ���B�>�
�r���ԅ���ݘ¼�0�w�v�p��m]�NV
D�W½�1�!��as�]H�V6@i�� �xg�����W�@΋�vQ�>��&�"���;{�_��x�� 9mG�JҎ�8��#XR�Rj/i�槎�?:��p�m�PQ�����S�c������*��O]�Wލ�k�܊��[H��y�*�6����|;��x��=j�U�!�{���C΂4��֘�s%�-�����w�z�m��?�_�1� ���1�Dz�YҚ�]g��A`ā���|�f�ΌO��vE�9��Јn�1c�P�c�}9�Xj�[�5nϛG�Z�qX�0eP�KL3�#�����Ρ���0�J�R���H�e�Zҙ��$�-/5�@D� �sL��)'s��_e�X��5���Р��,ɂD�J�:Q����co�_k��F�����_ �&L˦M����{PW���!�x���g.����k�Y���p��@+����$a�,}�byIΫ�IE�;�&x�sk�rJױ,3SؑA���ш�Qd�w�r��Up��s��%���to3V1Ծ�G�zR׆� �l�k<5��
QJ�s�͑c�)Wԍz�-wsk0��#�)Ú�S�ʖ�Yȼ߉B��_�GX&ˤ>��9�GA᱁�
�h���#��$A�y �>�=g��_��4.hU<�<p29��x���d���4�������¬�5�Ϻ�q�C�HY锜gp�,Ŗ�,��x�8��ԑuI��F��h+��δo�%�/�xH�f�8sr�����m'P�"=���N5�Kɻ��c,���'I�W�Z�@^�حJ����*����3�E�
�<�$�L�	�m[C��O����`�E�R��a9�m�\s�\�G�T���@Uݼ�p6R�4��O�a/�S¡&H�z%��ۥߟ�9�p +�8���7^��a���n/<դ4^A�ɛ,�o:�? �S�"�ٷٽu5��Vo��O�-w>hg�:�RID�x��;f���]�+�P��ߴ�|)A�x�3ƝQr>�����jO,<f'�C�[S�#����T̃a�.����� qp��.��G��$�"E�ܠ@G�D�rH��A�f̭n��4���3�ˣ��ǹ��z�4y�f�N���F��=������0}�����`�B�s���E����NW/�I`�A;L�AA�w�0�������t�MJ#���4���e�A���f��.w?�:-�!4 8�/���͈�Xu�T�"2!`�B�ّf�#��}�{��T�CJ�7�{�͞�Qo#A�hC�;��vQ#y��BR�qm,˦־��z�ȝ�|ABe��ZGoȚj2N�;Č\��w L<�`��	W���s^���Y"b�:wҺ�\�	�)Me���~=�:������F��>h_3#���,<��ؙB2^�����/#��O��/�^MO��< {���B�M����]Ct��Y��CG"m�0[�(�O���,.�Җ���/��*���^����/��G&4�Q�
Oҫ�U쪺��oS��!Pv7芋+�L7ca�6w�42����e���z���c�+w��QA�w�j�#��q��7��k�*��_	��ا\�.B��)c��/kq�����hM�,�p�(��K��u7�m��N�m�9�~Vr�&V�7��V)�S�hp������e�:H�*�$$B���Y�����F�P|(al���cn�k���p<D���8���V9U̺�Po�%��3��K/���Z�(���2�~�>x0�%1��H�)
���h���d�4@j���}�.�39�?�8��hq#$q���v��F�[�z�2�9����D:�pj�#M)*��Km#��d�j��\�v�s<�Ҭ�$���7�&Ŧ��p*�Em���3
�c���~����)��ֹ�������s� =�d���N������P�E1�/#xB�=�Q=�>�@CW�;a��JX Y5��67�/0ւS�2%(h���uZ據���3$}�knF�B���@���]�QS�ų8&P��\�}9�� ��Y�͓�A�	+���_2�>��A��UɃ�G^<P���?Vn�!ג�����-���注�E�s:�?W�,�S�7�Ԛ�y@�%O�t���ep$��-��?��h�S ��Iy���d�Hu˫�������e�������+9��G)A��0И����ӟ�N�+��"�9��c��'V��ݶ���!�8��{�u�i�5V*�M�߸x=�:^~
~Jۣ_�"��,K�g)ر�s�݂�����V��OT��'�;:�|#į˓�VwcG_ƫ�P�Hڹ%n.�+���u��S�+3>�W=��\�n.V��X�Yo�[��hdk/�El[{	Gʣ"�X�����R�������C��}B�TCYa��i�*�W|��j�����cYz ��(��A.~a��r�~5H3R�j��"��^d�$Z�=lX�x���(>Ψq�guϩ���\��7�ܕ�g4eئ�e|���I�i4KH����d��d��H�KP+V���^�qr�Vi�Jo���h��Լ/�a�������pxB��ڸ� �&8��Ӽb|�<��&\�X�.�g��+���EJ����ְ>y2煃��w��gO74�i� "�7�0�B���I�FG�ɒ�]�VB�$��@�fTمD�����p�8C��uK�O������'AtE2�'�j?)R��8�'n�e��.|F�l�L��u�{(���p��\8-\�;��>b��� ��[���W$���.�ɀg��N޴��$�C��IKe�#j$6��7�(�e!��3�k����F�C�R�#��5����߳�"/*ۿ�ｹ�������PM��	��5�Dc? H{�E���'KوZJ�G����S迕����������P��֐��d��"P����i��Ϊ:��R:�jq�Y'�%8��8W�Vu�eσ�/Ą[��[�D$\��Ç�H�2j�C$��w!�����2��ق�S�O#��H�-X-�����|�ar�^`M��c�Y�8�I����{!��� hֺ-��ۥ��f��R7���<��׫f)pT-�B%�r���	�#�en컭Glu��[�V��"��S�x���)��-!9ٰ9�y?�סC&�N�|�J͹���c�>J5�@f��b7��L��e��~h���v���,ld���Ot�v�H�p��s���b�f��)������&�錩Л����(9�0�vZ�c�]�����5���k!��Xx:c�W���2�[�4y�Y�^г#"�^��d�R�H��s��lA"����4�O�u�:S���lYӓ�{�n��n��	��2F%sڀ�{�#eA������5�J�ϨM�\�� 4'R��.�:�e�#��4�ӢfjcN*�������t}L@GHI�r����~���s:#"��6�1ilǛ�s�\Zm�%ӎ��ط!��U���t�e��Dkc&EOE�G^�tVa*h��B�����j��?KY>���[��Iȴ��[LC �ϰ��v0&��'\ښ4���5�[-ظ��G)n��&[a�"�ne���N��U�/���~� H2LY>�Z���q���M��b�.����t���sn�6?fUV~�54�pr8���Q�d������K.�\�e�/�͛���SM�x~�	9(*jk��e	޹�d1�X/Д�A8bέ&���D�Ý�ߋ��-�5�~vǻ�Mg+��#�?���?�1����H[�ba�'A�x�+�JO� 9��qh�.<�!�@���n�
�t��G���7u�-MH���!���ou���k˧�
�0R�v��=><�s���g$3j�"�x|��Y��x3�GL�������֝�����e�./ĸ�yyR��A\�8�υ�k=����~�n��=)^C<�MQs
G:�<-_�L�Z���H��y~�Ee	�I>���]�#��z��^�{�*�6I�HE_���;4zJ;w�`�*s���g�jy��:|W!'L��G1�@T��TA�K"{H��T�Q}�Y�����T׷��m	�I5��}���G`�}yJ�^���p7����^��[I�C�D�����U$�]���b6��Ą��o��x&��1<��C��[���T��~_�h��<�f��ț�X�k}�GY�����o`�Ĝ�ϫ�P�E*N����G{Gk�H��M�]\�f���`=�m�S*G��7-����o+�meY�gA�Q�C�/�q.���YaQB<>$�c�o�the>e�[�i�AYΪk�`w2v4�㫠�k��x��i^6ǔ	(n����ԡ��z�V���]=�Wr�^"̗[��ts/�2ӭFC+��W����m�D�P�gw���"㛲({�4�J-��U�b<!)�b�p�O��T%��i%5bA7��^B�%���WJ�j d�A����}{bJ����f�f�W�	�V�V�y�O�p���w�6��oM{m�j�%1�V�<9$ev���)t��Y۪�t.�&�ǅ"�n�Za�)�(�y��RIy#�}�2��7ID�q�H��a���H�~�����5O�,�.7�2�ĸ��vI�\��N��T}��*�^�]B�^x�U'�ۢ��7�O�8���ҥ����i;�
�W��m��;-p��Re�d4cm`�3�f�����g�4}�'��|���l����,Յ)�*�����7�k����/?w�S}eῥ@��{!D��?�1�O��(�`��/-_�[�l�}�$�n���).{Λpd�a�B:��z��TL�G�9������O޵���~wj��r���$P��5�%�㾤���(�4ji՞%,��Q��8���䶯�����U�v�B2x �z�y&0F�3K@�ȩ/$�k��8@Nkz�A5,�-a��4��(���_�� ���d�*�ؽ덦8���`C/ ��*%�K��D2�op�;hV4N|O�®�V�U��r��O�|��J]OH/g)���w�loB~�퍎�Yc���m������H��|��%"˿�2ß��X���`�4��/J�x�:o(�X�nҗ��ݟ�z��#~��ănK�)���3<#�V�]��c&�qm���G����'�e����{Y�v�zB����q*������D��Bae(�\� Ғ�	��EiIv�
n�fj�zv�!	��ϕ���s:�L��.1�l�f��������Cq�n�i-r�`�����m���)����G�ٽ�
7M��B�$Rp9J�Q�r��R�}�JO)sU0�rͥ�ȋ�P$gmp����Q�oG��C@�}�������:�}CwdI��%g�X��`��[Wr-���_Q���@��~i9����״{MsyA[�zG�4J��=6$O���,�[3}�N�Zm��/l�ŋ��Ӱ�Ԇu��
V �x1�ps����s�93.�F�@�`ٟ��(�u�W[L����x��V���[R���-QՋl����ϟ�h��-�h���?���.%�j<Վ����!OmcP�2cdB���:��9��(å=Bi֦�k�t|��.�����1��I�m����t��Py��ՄD)�-Yj�	�kҥ{�<P��ƫqG��R���nC��ӷ%��&��Cs�~��<��.����6���4}���&������f8&����x��r 	�,O�0{H��gP�{!I��X:�g����U/�T��E��U(T�e
��kNg�r��jiI�w*b��1{���tf�|Nؿ63*�2`�B�_�.�9>Z�Ǽ�7���^�YE��������M�A��>jB���N��H|�JwY�P��8'���_�]k��J��.���ȠR���N�,��HUҁ]"��+������]5lc�A8�8~0�Q.t���.*i��'}�eRZ�<�ʯεQ�A�t�N���mQs�A��eϓwg!�Tz�Pe
CKQ�S@�=���u�N
�"��Kn�4e)��>��YG���u4�݈�1�2D�/�0ӱ+'0�$�(��Jv�A��:��`*@vxW^ﭽ�V�i�<r��P2��Ƅ6f�����,��x�^�p�74��dK��:]�V��'�����K���Ћ,�E�}�X.+�d����a�^�p��N�b���⹛T������)���5�E
�څzP0V�k����rk�5���Q��w��Q�����i�am�V�:����!y�3WA��̓�yo�4�\�X8>���䈔fY�Y�q����!���iF�͸��?�I�z�2y�7}�P�ߝ\\�Y�f�([I��l<�Cs U�X^/@Ĝ�� ��Vo&�BN��h`C�?��U�,k�X*IQE�e��{Fn��)�y�M���a3zv�e@t����y
q�ތ	^yIyR�:�(�ɨ˔;�ii﫺��%3�Y@��P����Y�D�OؗT0�o�>�D��t�\�$���r�M��g�nQ�Z\� ����}�[���@t�&�K�В����A�ۧ��_L�b�6�]���\Rd��«`�&���ʶj���o���B_�D�������a�7aK�%m����#�ԡ�:���=88(G�X7��*�7<�H�����_먍O��֕��@?_!�g�vZ"\C���
��M3���8�#⮶s l즆��F�fD4�#F���^����ۗ쪩��{���n�7�����\:Z_�Լpe/��	���+8�C�K2�nj�{ Y{`ZX.ν�g=����U�	�dR�)�� U�7Z�1���rz�p@=IM^˝���%������d>�JU63��x3�+z
�_���y�^%)��3k�-�l���H��"��-���OסI?�;cQ<��T�1��m7�XVM.72�1k�򏖯}��.���0D��^�y2��K�.s(z��,k<~^�^�0����a�/�R�qM)��H�rnҵ)�������5�N�ne��(�7"K�d�F�N�U�d}l������oՍo�$a���t���4�l���|�ޏ%JĊ��gNV�}�&�S��js�#%٩=�$�M�����ŷѾ�lm�ϗ�)�f�֞���+zM��a��r(t�"8��l�JFM.=�������b0-�SD�~~Wn;R�0��O]��sĥ���Ŏ7��(����� �H�D����OAK��t�$�/�c,Qh���aj���q�!�mF�������B�|Q6����j����q���29d__�l��Pa$`|�xn�"�*����T]v)	����4݈w�I�8��]e�Q�J�aC'�j�Ql��0������I���*J=ɶґԐO��&_J=���*U���qP^CC�Z�2.Dcԡ�&��>-�Zi���oq�kc��*��k�V}b�.�bS'����m�fБJ�&���=�������'�?�Wp��il�|��E,�#ͪ^��iN��_�ʇ�y��.L��4
6 �8����4����0�d�C��N�0��0�J�'�r���_�A@���).�:V�R�(�#�rܿ����0-Ѻ�s~Tm͔��m�X:�b;S����{p�'�ULa�ՓцRgbt_[�ke=����޵�Q��d�yɛ��7���%xq��b�����f̢�r	5N��V3SJ�X�^�+��@�P�%GX�P�}�g�.a!M4��B|l'�/�ޔf�Ѐd�����(�q}��pkMf$ov+��U��3A���;٤Jo�����/Z����u�UN�`�O�I9ֵ[?	ZZ�aE	.���!4P���	"��rt��?6n|8�4)��v�����}�	�*-8N4�3��e�K��g��ud���kz<�~�B�*��/�̕�a$�d��G��e:��
D��wj	sEȍ1J�Y�Da�K�̈Qp.r��YHM _4�9Ϟ�r+��_�VDl���a�nيx�7�}�A��b�䲟1�#��D4Tc_�ޥLթ����Ʒf`��H�JO؊�ꥏw�w����l����n}$�#ܸ�E[�ԏ�Q����JN�G�2�O�X�����oo�%��w�Nh����]y�S{VH�VNj?���4T}2�9v:_�����&���	�7DZ�3�\'睉�r�X����a�[Z�̓������Uc"�4�#�0Ua��XX�9�5��Ϝ��?�^
���F��Y4͆��ҵk:5�7w=.���/K�Yt�E�hE�*��)����I�EP���P!y�ᬪ;Te릖���PZ(u�qؚ;�hyn���$�Op�v�'��9go��E�q�S>۫����}ח���>��U���n6�6�H}[t��|���=t�çz������R�)��L&B�=��Ϫ��j���µ�r+������8�n�����i�����P��ML��� 51n�?���fx�Q���jY*�;2f���j5&)�s�ק���67)宮6���վ��>ă�~$ۿM�wvwIG2Q��k�g����|��ԩb��lu������ Ȫ����F�	of�3�a2:�4^c�#�y#d�F8��X��(2�>�[4qm�ڴ@�+
�c�1��:B�r�a��^q��p�X��X����M�$�ε��]V��8#�	RR:p��r=
II�PW� Y6��$gmæ��9�_A�
�?s������F�`X5<�;�2R.�O�Jy�hO�D���h��Z$S�l�\��$ �I���"��K�8f�`��Zv�
4��Ʋ���YBi�4��n�a�Y\{Y�Υʧ-q�2/'��U�0(����s�50����hѝm� ��Gj�]��hj��D,�k��l�)��Zlnm�L���9���x.g	�|��s��Z�{k�}qM�D�6�$3�F��3�q���w���K�q0����Zr��
�E'�p%�|��0z����������h>&�	���J�XV:��f*T��<�bwD��A\3���,�<���S�Fn�gCW'CC\����)֓Wʗ���S�#���BK�ė�c�}&���)����o�x�Tu�T��(<}�2�6�6d~̴"A���d�귘t���+�N���ꇧ���C{V����m��.|�ޡcXۃq|l�H��SM�n�n�=�����Hrj��B����󲀝i��,܂���<��F����8�]C1w�Z����29Fj��r$O7�
�S�龗[���/{7A� #;���bRG����t����"�P�(=���z���;=��v�_0���S�΂�7�9qi�eo��3���$��f+��7�:n���;*��6�� k��Z��i��՜`g�� C�AN���Ja�Yq������S6T���������kۚF�� !>0���������|P���uw��`���.捂}%.��>e��ݧ+�TjR�}�f6)��3�7ҷ���߇�P�&��Pp�9]>���=�z�t��r�Ɍ��@�ײ�O��V�m�j���w%���_F���/�yD��4d��;=��菏M�_5�w�1ҙl�
���fu��fo;����+���&g����'�T _F4�ڧ��݋Ֆ��9��2�ļ�>�{�H���+���+rH�)��	+��*:|��gb�����n�
��Y��њU�5�M��,U_���:2N��fe\L5�qm+9�����.����C�.�b�Hf� ����;�%����8�'ZS�LÃZ�/F"�����i�nNy8�4��z�sky'�Ǿɫ!���"�Crغ�N�(Xr9w�Σ���P͙����Ż^�����w(]��5��D�+�PV�ur�r�RX��n���z86�����K�S�[���}nY�x�[�~�y�/u�Q-2�k���Q��=��c�v����c���,��*6Y��U&|�I&�+8��%�/,��Ž��j�us�xn����ߴ�S���:�wt��幀m�p�g#�iK1c�<4���/���F�e$��y}2#����/���[��d���,��1�ZUo�;�۞y}<��'�?Z�S�0[�y���='�P���*���U�p�s�C!hS�	����Ӯe�q��U��^��,��H�F�9Z4�KP��h��g
� �������A��c���f�1=��>�׽�x�5��g:�����=��"�D ���pjq�Ay�6Ў^�7��ϪE&ˠf�6��=ز�m�o�sjYq��� �����p�p�1
�(���ZS&jj-ö�<XHr\h$���RS�I�|��U!���'����H�"�����^;ڙ٭a9��pnL	;���8�C}�;�
1����yrَ��]v��Bi���!��w/{[�ś�:Nz���F{"�er��K�g4�%������?�Y��2�r���X�\�I����@�ӄ��Oȣ�Ik��dT�t��MqevbA�s~�h��k9�Juٮ�T�Z��`}8�NA�H�B�5���¶y	27[EFFM`*u/���y�1#��&6=�o%Vq�J^#�Gp�wR��(�1�%*u~L�D$fe�����*�Te4߃�OE]XK*?DVy@�R10�Z;@�_�!tp^��}�Y���D{��0Ё�F���� .2�;,t�őG����p�{q�d����b�����<�_L4f��ڂm~'�<�k3||��+��,����&���a
q;܁�V��'�r�9����	N[�V��S�yz�e�b	��WQ�� '��i��J�B|��i�$�D�/aD�2O��ծXY����[@nߺW�R�L��l���滇�M�V���|b�٬&����
4"xq��TD�r�����8�+k~x�#�9ĹZ�C�[}��:j<T-#��h��)(�ӊ���O�l�^�a�]����Qe�K��:��l�u�Ŀ��T�^�06֥ K�%*�#�?
](!՘*���6D��\E��T7�_�9�3`G��C�3RwC!,�I�)Kt"�$�K/ꔧ�`��$�DV�q�6�0(�~�}:g0h���5�lWt`���>��(�21�W�����d��%QD�2LjL#��X�.l�R?b��H�zW�(!Hqd�=�BTa�qg~�p� ���5<�(|F�g��)�l/�4II%�g��b�>��"x��Ӱr�Oq���x^ׅ46�8g��3����6(���cF�L�;���Jƕvi�(��l�n��8^��tx�̇HK1�2��V�����|�8�p*�K���(����trJN�P�!�ڿ$p,%����'��xF O��U �R�����7�^֗8RC=��$`��]8��0��T��C�Y���v���;.��(���X�iS�C��� Av��F�	����s*I�>Mm�����I6��0y}�����Vq�'��#"ߡ�R��0:Nxr�϶�'�j�����_�U,��K�+�Q�9+x�:	�-F�5��OCۣ�o���f�q��"�f��C�KM^�0TȔq�)��4I��f�3���Q�Y;rq7�����{�wUf��3�>4x����?Ir���ڋ|^4o�����@�~�d�̭L�]�C�v 1�ή����2�V&fw5��˂�E���-�G����[!l�p\�j�?�L��k�Y�Uq3�*�m���@Oc°StI z�ۓ��{���9��;���{"�HG3��*�Jq]�W�%CgZ*2މAQdQ%��~��Bt�m_U)R�"�2ev �UvL��n�z��r�1G�����CQٝt�'��e��HT�N�dr �^�-~-".��_�)>�hkY2G
4�ܩƚ�L��%w��/�}�l	���B�K���-����J�ˈu��_<K �O$8Q_� (�l��䰕�qm�m��F�N���lJ���X�
^�:t�����+�u��㺳&�/��o�w6�b2�B7W���Q�hy��y$�d�v�&�<�Z\���7�C_��Y�����z�s�`��.�m��讉�}�!%�

Hw��4�{l.��y�k���5M��� �p_i�zpdjbN��䯑�=�Xh�¬��1l�ً{^T�������-Q��K��H�<OKP�z�GJ%��T�#;��4.9��~�N�g�%YB_1��7!����F,����&f!�<?8��q��o襍�C1�v�\�PfN�m�t�;�܄@G�!�B��I�O�;"a�i[�X������z�{�z%����r�����:���nl}ǭ�gf	�r!đ����	U� IW1���&��S�m&6��ҁ�T�D�y\�ɶ5�ē����1/;��U�&D�����Q�n�7;c+�<��k�ֻ����o=@/�A"�̆.ţ��LF�-M�W	�n:�	���(L�;I�w��oʽ�tIM�e>�t�t.dH����پr�!���I��B~V����>uf�r�q�
�9�}���eUH��Q��xS�G6��/P)����J�>ڈ��ȷ��̺���L���X!E��N�p�v�RWM�h���x�I�89iD�^�c���U��y���o�s��=*�WWM�92j}�u\�i g��c��y��n�Vi�O4;��ws�:I$�e s
k[8�~1��n�n�KC�㢑S���~�W�r5��N��ǈ�:�l����Heَ�Wl����-G��N�:*����4&`��;��%Ԑ,V�,La��3�ŏCR��z�0����������{��ŋw����a8�М2�����`>��L�e8�QL��Q�
�1��������{�m)�G�d��I��svշ6�猂0 
)ի����>(\q�VnP�\$˪��z��Ǣ���}�[~�"kwRE�y{@{X��>8��q��K�&:D!K�1f����_k��ښZ�Z3H,���Tp����R�h��w�nG�jJGa�����lo
B*};�U���S�nW���3��8�N��z�a�<s�-e�5׾�����=�{#��$��}��CTC���zY��tTsT`]��V��9;�W�i_Mm���;��{�H���](lq�v�����W\Zfچj�&�u���m����6�z�R�ŉ-���ո�M����= w��^�{l���MD�8\�
��>�c4������\	������_����S�&��\����D�L߆U��#��	ھ�O	��M�;��7X�v��:�	�8$$����2V������=(�9C��s�o*i��*�S*�h�Z�}��d7�X��<
V#����*���rxN;���t��>pAM��^�T���Ē��&+̊4�mQ)8���uKf�߽X<ER�lT=��ņ��-B��/`���<�U���!r�
�=��g�'"V�J�܉_70����]:�?XUEW������7�p?����p#��3�;^y�U�bB������$��HI���i�)2V�5����-/=O,&R&I<^Ʉ:�ګ����F|A����lF|�]p`D';|�H ��)ˣϟ3��~T�ŗ��{��%�yBl$���$��s@Ԥ%�XJ��{�$��Um�~�����e��}���NP����Irg����)R*��?�x֭J�E�xx�2ҕA�6@��A���N��n�
���[f����m�V61�����^�̀�ݎ��ە��u�Wz��ѩN����j �XR7�dÏY�Y͠s$���`�88M@�*�qcSx�3\(��<��l6J�n+U�c8d���`#�Xu�e��0|���jίh���,�z�0�M��t$��*Bɳ.�W�~�_��_�y�&��C�$�b+D�;�T�=DQ�C��RR(~2�:��V/�=�M6ti>4J99b=;��Ä��N�D������<V�k��� � �H�r��ךlw/���@�4yp��#�����W�B��	�m~�d�m ���~KN�Ftz���\��Q ]�����f�}��*�l�h��BRlᨫ�p����F�P_';��EO(Gl9kc�P�o�o�����O����u���3r�{]��i�*��=MV3f�����v��8>R4�Ԩ��4��>��p#4��Ɨd��H�G<����7���� 2{�̓�Š ��Qk/��1W�����K)h���4(���o��"�{��?�,S���3�	*"ľ���{�GiEU s�_3�	!�(E�=���ci���nb(��o�_��a�c�b����O�����T���ҭ�V����	���
�*8ǩ��S��4#S%<3���rs; ���r]8J�E����&(|;dh�a~�F>���B��*@Ķm�ڷ�����_��{L~X;�2�Yq��,�#T�u|z'�W�U����<2�w�`X��� ��� ���]��;6K@^��;Eș˶~�P���-慳i_���7_s��L���d䨼��})Y�봴M0� �!>�NP�Z?����ȽꞐ�׿bb|\�݄�Z�,��9g��j��>�,_�4�����b���C;�y�t����t!w�lu�Y;QJ�v(����_�$ڮ���}61r�h����~�%	D
;J����P\��~��2 �M��
��=F!������\�-��M�9GȈ� �^�)��c��u�c�BΉ�-+��*��s_�t��~�+G��l��
�Qz��;Yp %���1�i�h��K+Á[n�V���ƻTv*@ �M�;���"�[�9�B.҇%@3*�\�5<b{x4T�U��HD������F0�z�*9=�m�Ƥk���V��9�oP���]w&槵ŝ�ޅ�Z�@��0��Pu*S�s.��hU��Q�h��C(r|��m�ہч�{DN���TM>x�d�ϟ�wO9L ��c��Q۸���th�����*��^�R�Fm����>�M��m�_��Y��@~��c����Z�	�#k�����:'b�ŀ;�r>C�ی�_�A��ʎ�Z�8sƼB1��� 7؜�|� �PmG��B�ߌ�QvY�9�c�7�C��6LLzR�y�z�1z���+Y�M�U����ҿ���İ�)h��4��_�L:� ��>���L�[wW4<���nQ��x���������Q6%�����+�t�� ��Ig��c Y�ݗy{�u��q�p�t�Ҿ8����ɼױ����`�,����^#�-I#zS�	���؝�q��m�4ɲh�X�}�ǯ���#���4d�@��8��������*�:<؜���"<��>����a�k�㗮R'�ńSS1񪃱{"�yx�j��N$Ji�T�n�:����p.��(�ŕ?mL��3"(y$���f��˖) ^����=�ȩ����7$5ʾ���������]�M�YP��mh��L�ύ�2P)/nG;�ֈ�VG��f[�(��+�R�!���`��$�l��H��2	��[nY�X{��;%K5�,?8	%���՘�I��'ز�JYI��Rj�����x�kf?Q�\n� �e���>F������|(���B���d���G��HZ��*oz6���F]~���՘֪a#���bf7'@BW}��:<I$����}�m���{A��~�-�ᎁ�Y��/�=Ƴ2B�b|��A|��h�+O�f!���۾��2�߷�?X�v[���H�v�wM��m��3�E�'���J�F�f���=+�c�d�LѮ�Rȇ1�:c%��s4���E�w�E�UV!�mLj�1n@A��}�2�lŸ�IC�B�T�nw���yC��h�8Fh>.�`*7jX�$!:,�	}u.��n�<��?�� 4�ȃ�F�8B�D���@�Z \�:�m�W�q��.ғ	炅z��bHi�@|�XI�np�\���u�N=�U�����iV�e���F�0� �o~9~@���?x-r���{����'�?E�`�͹JJ� v.}�@A9�[=e�k��q6̅Om��.Y�f����1�U��_�)�+L��a�4Ԅ�������I{\#h�$�0����s�'.|&�E�s�/QK��h���i������V#8�tB0"�����?��׃�%�>�1~��s�s�F��������md%{�Y�,��Í[q�I%�e�`"^�*�%�`����3�h[w�� ��UO�]G���(~O	btYu\��&�P�0�e���-�����}��'a[�/��V�J	��l�G�g>�O�F[&mFn���s*�x*ǎ�2WXL_@�-Wpdؾ�o���̷w.N���;�y�]��+�+�J��눆8�_�7�OA����Ke����>�F
׿'0�?]w~ޛ��+i���oƂS�}��n�h�"��n����$��
������g�ٶ��xk���{<�7�⑅�:`��E�3��r��R����~s��0��ꙶ�P�T�ikQS���@�I��������\a�,����䗒��:���g��#��vL�u3kTԉ[���Ftʭ��G;i�N MC%�j�����}C�B�5̑�fԧ���B�u����?�;7�Ք�}~�+a�c�^J"q�g�:���z!Y�nNQ�B ��CL����|>�Ak�C�҅��+�Rc!w`35C�rv���{����wn�V� 2�G|�t�ͺ&�1['5�e/�[1�!��>�Dg������2m�'mя�����G�����l�
�&���iDngY�nr\&D����+_�>rb"R�͐vui
�K
f՗�k�o���C3LRrz{���q+Z{7*B�OZ������MFP�?/�EO٫����բ���]��:��>�k�I��s� �Y^@	�*��#��,R
UH�ʟ��̪�����w[�6��`��X�12()ff�>%X���-���W]*��g���N�	��>%o�	��|�,��/�������/��C&Q��=N=�N�����Sh��T��hz(�������JZF�\�����nE;�[p�
�qb%Lg�[$��V��^5i$q�T�0vX#�u�Ĉ�Z|�{�(��������q0=Q������0�Rچ�Y��y�Kop:�K�#Mh��*`��'JT���pw�����P�e% t��v���휡��� �mb�&��t�a!��z�/�q"j�V�w�dn�`J�[lL���Ab�wN)��v��2l}�Yi�e3 ��M`�T�$�`����s�ʚ�� �<���p�Q�����XF/	r�)�O��������'@��}�Ü�S�/,�U�ط	���X�@T�t��a9Tn��E�¬�U�5<�V�k����9lr�tU*��C�J�h�iO;�Ȋ $̦��5s�)|�*�1���xAuG�w5���5<������!�� GN�l�q����A)��e�lB~���^U�O�@�ؾ��$��W{��A�|���Q�����M8�5X�%�E�>����7�9�N�����4�=kq��e��>�/��f��>(�5𯞉f��cm!bD�>���J{�:�JöSS������n�D��V�vAò����m4W�[?U����>�v�P���ϖBs�Ղ���V�����Ka��y�צ����V�ٿ�\y	�z�8CĘDiW��J{��$Ъ�� k)��;�������a��?N���k��F�4�'��-W�uqwR����`��6��y���
�l��4�h�W�:�Q?���N I4�]0�Y��	Ȍ�UoE7�q��c�=(��TsD!�'�x�ŧ�p�\W����H;P.<�x�I/;k�ʤ�+IYME�^�~K���(j���g-�h�֨e�,���āW~b��U)��a�8X��w���B�a��Jef7{a	K���9@S�����5����/�����Z�0/M8��N���_�m���(�$4����he���7�f$V�/�M���y�����vҡI���T���
6�شP�N����	e�f�|O@�"g��E�g䆼�Cn�J�j�ᬓ�\�h"��8�PvZiC��;�������8�SG��(�5��/3�W,k���N¾�譐N���Y���,��x��Tm9����5r⊁P��3�W3� 3kz�,�����|�k�h�%񧮴]a�M�d�U���εo�'�N��ƻ%,���l(�9I� �o����RK�3���ʲ2MEo��5 $;In�{�F�S�&N=�r�" zD��N�(�	��Gw��JTe�yo��:n�L����f#��3W3Z��7��b �j��?��@;�!]��D�\�h\sנ�+��խ�����"��Z
���V�tq�Dq:9�N�ݘ�vT�-��^:Z̓8A��OD��d����u-�&x!\�����d�U�|�h����K�\EJ�3%!��M��?&�!�@�v���P�(!t�%Oc�������>�g��C �d4���w��R=
Y��΢{������ձ,n~��\���~�7{pJ~7Qt�؜޿[�=?���l �F.[Xۭ��d�䄄��vpw6�S�_�od�P/�qy x�Y�N��⥦�JB���I�;-�d�Y���Lr��4u�<�!o:.���߃�fH�|v�/����A��`��Gl/r	ѯ�7\���Vv�6��Ϙ�<!g�D~�l.�/�TSA��nOQ�M��ͧK\i#J���7q�7��\)���;���>��J�?����F��|�1��{��J\ �u8�s��))Wצ�u�;�w�o	L#ϛ�?7�Œ���)�v��{�;�N"N�i�j_ %�[ڨ=��C�]R6�x
��hV�O�i��G���}B����"�rP���Q?�7�(���̲p>\J5bI�!R:�~��p�	"}������))��I9i�_g���%
f��	[}hR>�IK�G�.�o�����|G��O���0I��P�6s�A����=̥nps/%vXq'�G��v�5�S�0"�b�,1�vf���Fde�W��׮">��ēl*�ZzbO��td�h_���i��vf���KXa,����-��C� ��� �y雘5�ͻDu�."��\+��OY������Q
y����{K+T�m��$VezhD���J�5�z<�)����"*4���S�j���"�k���,)0YQ�
]q������n��AN�6�C� |�z�J��C�ǮU�����4�����KL��TCΉ�
I�8(nĳ� �ئ��>�\�1�%�UA�v��Mc@����H�+O���[qqD�g�Ys��/���/��yq���VYʌ�@?�~�
R�o%�!p28�[����~���bJ�,�M�p6���=��\��q;�*]`V/Q!�̊��6��G��x-�TU���	p����1���zO��H��Wf��(|���8��2n��	3�/�G���τ�v�"�1��oj��Hj��N�:&^�,u�~T�0q?�{��Ә����/]�pw$+�5r]Y���ק�XC��D�J��.iw��
��[�غ=-H<�0H	��&c�콢�> jd�!D��¼��rY��$�Vy� Q hE݉E����}A�\�J��c큈��S0G���PL��_��⛡LC��灅�|82�n�h
JQ��ee���ν4^Gf��9�{��]l��tW-|4���o{�%*���x�7�x�J8 ie���=8$��f�~�TT�L�0a�����^�1���`��մ�[UVgŤ��^�I/���Ƒ�A� ��%B���F�q�AS6f�)�����V̎�i{�ؓ�k G/�����@�ˏ�&o�qE�i�­��ŹK�4�LH+��-��Q爳@����9m�2�a��܍f����;y�,M�2-�Е���4EC�SCh��u�PG�Aj�<���g4�P�x�G,������f��C?���P%C���jFo�ܳE�4����0�&bo=\BRcgP�q&������t�Z�S��uߏ���.�&���̨���
�!�
b��Ж��*�r5� [J���|��Md
�m+�"#���":�\��#n!��q ��������J��f/�t(|@@NrO?ݷ�hl��[-�Kc"P�CPXh�bJ*3��^9:��TZ��0f9e餛&$ZB������7�����'�L�T�'�!$ul�9<���[:G�*�j�f����Z�ze.>�DU�v�s��I���}M���K��l(
��S��/��}��w��t>�?����+ {����Oi%���s	��-�oo�Ǎ�3/~5h���%��?�/e93�1u5����V,�;�ձ�^�SZd�|���&܍�w��	� ���ꝃi��B�
r�>����.�ms��;�v�>������`�
�����d��a5�$q��'e?����\�3��"�p�5�ɢ��QT���Ws5|�2� ~�<��� ��\ҡ4ܢ�D��믴{톏5��?e��x�NIo_�c0�ܵR~�ű��t��tW|u��NXq��%��EW�A���(��;e	^��=�B� 0�j���	m}X#�Px����uV���Dc%ӁF]]��A4k�.B�ш+@�x=o~G��m+WAh
&-�X�u��A��J���J�^�fԖ��I�o�� �̱��H���m{i=x9��4��CT�ZڣA\9��`�)�Q��:ʇ���h�*�=!���h3j��G���Аo-`�5j�G��[�T/>��������O�Z]a��q�?I�u�F?_wC�DhS,b�5J9I)���O��$���q�X�h��V�[9)�VF��+�$I����ՇG]H�~Z`?�g$�40�e��|����KWk�h�+Ug��-9I����b�JA RI,�'˵� �{nq�g�qufl7�%����%�J�<���4���[�Y;��S���i��:�L��.�/��9�����|,��V3;�<Z�vv<(UQp�ތ�݀X���lj0�z����Da�+yS��H���oi�Q#(�px��!�����[J���1��9h�ǅp�&��X���{�a)4�� @�o��RJ $1Q���=�����_�|���o'ϒ�1�f��� ~�@���A�w:��'������ѶnmW�%{�@q�D�F��P�8�nS%����&��
Y����
!�����~�$�K)Wђ�VP�3�ܘC�tF��qZ��+�kC��0��j��l�����Mޜ ;��e�ʨ��@�������X7�aLD������;�Q�	��D�3��DRI���+>m�߄	ޏ^���`��a�{G{��L�g7�����^{
�g��	�ڝ�_o��n%ūG�!���e�E�8,��RZ��-_��DH���S����K��m�)_ ��%�zf;7����F��epK��wX�v@�����N!)�q��w�=`�e|���񇜡��PO�A��x��i�[s��a��)��0�kz�O�2zFՑϤ�g�'����.�aL}�&o_��!��9�h�)���t�2���kR
u���!�w��r �tݓv����}�4Y��W%E�ȅ$�����bv*��h������!�y��/�����(��1xJ5a��6q���z~cɃ�Z����$�f,��9�z���i��^��EBC00���^$��e�v�;Q;�c�\*5-����ykP­*�r��a $&ȁ��և��y�]`u�q��J��ؔQ^�;���
�-�Y��eMf������}�ȍ#3�	��,u�Z�&�t����ϫ�AB��K��Z:j����Xy]{�����D��"��w�|%��;�6k�)�֔a��	/o�l���˿�Y}�����I�����@I=0|�ϓ\F`"�K�=.�5r�(��^ldh!-��.4����Flk~�~iBsdwrO\�b�߬ovy��.x��7����%�sCU���WX'��=��
U�d��1s����vr�|�*H[��N�Yͅu2)}�5	j�<ַ�;����=�BG�'ρ�Z�3�ذ7�<��c_�bq�}������!�K�� <Vm
���f$K�0A�~��x���J��\y��s'd�0�V��iu�5u�B½�x�����y�Ē�]	-}�<�|���lO T�m~�:�XU	�8��)���k�Y�'Go��I�AS�6m�"Y�.�P�R�^t��Vy�����m��:FN�.�/�C����A���*�x�J�	Q��Ї�q�`��}0���,O�������h�y�*O�����5b&�"��-��>��q���Wf#��S��i��Z4H��됇�@HfT�ӕL9��~�A�_�`��N}`�������	R�L9j��DR��t��wokx�.ZKZڅ�	�XD�����h�]m/�0�<�eH�D��{1ᜉ6p��I���[`Z��:����Ȳp�>��fE�J㆝_#��ld�?�����0l�ۥw�Sٮ�m�vJnp{@,.�ဉ�rql�*`��?Z�o�>����8�XE.�ݰ���J��e^�^^C�EY�M�]�1N�G��B_���t[a�;���1�l��9Pd��H�g�!Ԡ�%��?C��|B=���^�d�z�x����y��~R	�������D�#q�=99��0"J���-�U=)�>��>~�������2�7a�$�����X�Bν<I��ΰ�l��F��K=�qS���9d�`A=���i 8k�/�	��Qb�^�π�!FEb�=�����T&��p�Io�9x/�����n3F��_��˥� ����HV�#�d`�V3��|�y"���XGdq��IjY�9�D�OBC��^%!�������J���ѷ:��9���m%/�h!A���1͐��v��'y }ʣ�[�|���O�G/��Ey��`liշ�yBq?,9Sn�0;�������j�[�1a�Q�+@�ʒ<ȥ1��L6��'bl�Di��|��b��X`C]��S�PC	/��ī�>"t��� fģ˖�<�����E7C��6�<�"�4�%{K)�\̼������k�׾��1�=����#BP|;:�_!��@�/��h^8L�����j}�����`��r}}p��C�Fiݗ=v4�;��Ν���.�Ź����m�}�V�_ɲm�����) �jAL��6��I��Y3�b�'<m��*g%��	����^_��m�&�_^����햙���'��9Ŵy[�����z}	:������b��z+9�V(;I��O�O�ݳT�����
KэMwn�*0�I�&���&c�?�$��A��Y�ۗ��ɬd�D����C��Y��j+�d�b���	�� B_��������-������3L��cKs���� `�/nӵ��+��������GHN}�U ��Y�E���p����+M�I��>�y�Q�%ý��wW�,�"���3c���)b�5T_�_n��;��X�"퀟��H��Cj�8͔�n*�����!2o\����R���50s�ڶ�G�~��A3X#���~	�`��>I'dZ�G�o
fߴ�=��9�h��H�}k����?x6�\,�l���=�́/�gF��T��I-��2Rob&��TboS-��c�|��P�.c�H���c��Z
͢ҩ����X��­�Q�Q�j��X�(GӤ���w06t�?@ ��E�[Է{/�)�`�B@S�!>Ļ\(52��j3G �k{�?��6�U+, é�Ѵ�$�Ffs}1���2�ӏ�h��SV���ED�A-z~��3^�f�d*
�e�ވ��V) 5)mD�U6`���8�x���$Y�����Z	v)��	��╏iݶ�b���,'܀D��v�˔.�c|���S�`g]о�W=Hc��?N��Wmde�Qlf�h�`ngx?�s<�v4 �=�!�*�I�auep��/�Jx��c�sw:�V�{�$o���i��n`����.h�V�I��I҄�C�e:��I���~xGr��پD�\�UW��/�L�y��Db�Hh������,I�F�8�LFP�_ۑ5]ʞ ��+�5�%��5��#��:�^{p�V���]��E~�ĳ�?���w�Y�3]�'��*����O0�ˮ�8�z'	Z���� )�e��[��v�/�D \ȓU� l(�3�(���m�h��eSu�0�]�
d���ג��SF���/(�a�ȷ�N�J�'�+ �ݐ���P�+�-��3.��Dg�+�0js��l-�~���>���r&�a{�P�Z1dh�ZR��<[6+q�P$��d�S��.���H_5%��`O&�����^i�ܒ����.�ϺD7���|��m�T���*�L��>(�6�!TलĐ{���G!���>�ك^�0�x��*�
� Z��Kb��#j.9p�?F4����.�&���|{��xv*}%B-=��ʔ��'A�q����|���6�0_��P�ۚ4��3�t��6=Ww�,W��e`�V[LmI�bV���O�Ǣ��JQ�����R^���d���G1 ��0�����b\p�\�^� ���](�3��s6��񮉜`�X_��2��tU�?4���U�֍4��Q;�T��,��K����	��-]&7y�M��7Q�i��%I��P���G ���֭��M���a��i���O�͔������A+*�@ӻKY��5�]WL��D<y�U�F��k��/'P��s[�W����="סa9�+N����O����/oQ}x $�dJ�Ѫ�Y�@s�yrZ����
���2�B��Jl B��;���T^��cς�M�f(8A>�\��!_�9<z��m|�ul�����܏����)R8�]]L�ФX��=�;B�l��|m��jX{A�]4X"�q0�r��:o��*�[�����oȅS��"�N��&|G�Jϛ�@_��/�'�e4�G%@W�y�S�j�?�$��^u�¡8������~!2MƧ��v�M&*����z_�H�Y�C��I���R`C+�rM�d.㹖v���ج :�|��y�Ѹ������j�2t��
Q�E�f�%�9���y���f-���zkQ�p�|i<��u��y�gfUͨ4�~76Z�V���)��k_�L��B��,��~���-km{�ʶ.�m���>�"�ă��KgkwbAY�&;��p��{����.>� 0�0h�QEO<, ����)Sj�(^y�>y�f2��c6���*��5H=%0�[k\d�2ڄ�9yH� AJt�6> ��u�)3���N�T���*�[�u����HM,��>Jݹ���5:@s�L�ޞ�؅�Q�9�+��m%巸��=���XA: �T�2�B��7�o�D�{b;o�u�J��ߵh+��4��EC��;@��/��3<�J��G�l�
��������srW�-I�}����Sq����'
�':�����u�G��s� �迖���7TiH�_q�Hz�҇y�㛞�b⧋��Q�E�õ�,((�͂��X[�¢��O���(�w�5P	�^-�����2��DJ���4Mު�8�o(U���h"0�6کg�(r��zj-���X��X*0��������I7���`�"����Fd��U
�_�;�!sF�%I-(�t�a�(��q�K�!Q��x�Ε�>�s�-��x�
ȟ=qA9�^/N�&��x��a�W�R��6u�F�̪_�אK���c�����](QD�x.�������31�k.��_��Q�
2��D}\XH60����`X���~�^ny|�%���'�:��d �C�V
��-H�6e�������b����w�ŷ���Si���{��X���g9���U�Q��GDiw8K�3����7.�b��_�X�$�H�P<89�2��	&����#j��3B_�� ��Nܵ�Éo���W����N،U��S���K�A�m���nc��
�.R���!g|KV�9Ȟ�&t��C�@wH�!j�6�7	gE����M����5L���[�;�'�<7�³Ν��J�!�6��9����G+
��Ŋ�*�Yx�+��yj ���Mw#���nDT>�T�5!�s8��(A��t>^���ty�ːѫ�͹<��-��p�~��cNQNy�~��M�2��仫�@�j���3�����XO��@1�v P�N��4}���c��nt��w�#h$[�ż�r�,���: ��ܳ��������U�>N��"FL%�E�5�(.����gل�����ZA5�&���v�'����?t�Uɒ�K����W�⟽�'������T�QUD�����丵�vbsg�)�O,5=�E�S���e��[o�9��� Y��Ij�s��S�v?K9�ڣ��A��hF�K��-�,���pQӸ��mA9կ�Br�Y[^��# �W�]�ˇ��˚��=�Nk��U/��3n<�GjRs���哈�h�BUL1^�j���E_<���2��FK�ߘ0GA�P�v4J$B,׽0���g�/�lG	s��@�a�����#���.�>d��<�l���r����$�Ǉ�Z�#����&S\��U�H�:����h۾Yo���8+4�A�N����JV&�Γm�C:�9�̓��`0�N|+��f3=82�&ݯ�M�V&QZ*LW���ih��<W���ĩn�QT4��������hi���Sv�z�?(����7T���w �-:e ��7|t�����frRK}�v��f�UQ
�3$��m_��� :~E
���N#��+������;�Zw�Ш0$� nr�vf��h�#�R'��홫L� m�G0��HT+��$���h���>y�+�����gy
DB����C�"���e�q=y����,��%��+��X+{5͖.� ��"�\��Cha��V�;�E��z���a��v�pH���R�4����Ծ`��ymK��Me�F��ߒ�4�4=�I-�9#�i�]�m�7��FMG\����ʘ|�������c0n��*�s�S���4�^��Ց���aw�@y��"�����U�mc�Dh��w�&���ǣ�� 1�wWO�������3��W?������˸�X���/�d���L�)�fu��NS�@@���1Q8Q4���t��3^���బU&>#�T���X����T�û�Gڳ�?}bƕ�mY�M�<��I�ң#�,�&�9��1�l�%��l�s�	�WXnT�>\�Im�-3��Qξq�%����T�f�7�����h����I{��)���J��ٲ�-ޚS�i=@�[t��.� *l*��P��ѹII�ktxкe�E�k�U�S8H.�_W���`����ǥ���Sopx�A+��9(�Fh"�c?0_~鵥!����r$B"��Y�x������R�&�"�B����$R�y
Ѐ�U���e�Rz�؎R-V�g�[|2ER�L���C���V4����q�l��{�E���ruՄbk�xA�v)2,D��m�
Y|u��C�NϾ��dS{e�r���0�D���}��%]�Q���a't����I�v�6�.x(�(þ|%�G�IDe/��"��n�S��jU_7; �	���=l���sOWB2sb��g�<t��<b����V�?$�yԾ�袻$/�*�杁�br�F��)�{=u���e!�m��d��1a� ������mk:r���@;�)9KU*�Bm���o��"� |��C��FҸ��$])t�\R	��@Ej�E���E�h�m�e<��gi���s� �;����?Fd|7��o�i%����m
Ҕ&���%e8��h��q��6���u·W.Y��kp|�$Z� G��ŉ2v���B�&���7W2I"��_,L�=��{��2��||#�Z|8�U ^���a=�>�*c�� w}��V�C�o�(��c�,�R�����2��������"�4(����}g����y�<�����bcv8 @�%�@��9j�̰��j*���yE4��e�,�K����h-YMnZ]`��2��O5�nd�w9}>��g���oS�E.�'��Q����g/�mƚ�`�}���B�+�@����J 9�ۋ{�hM��'���7�֙��/fZ�֕o?���vVbZ�N?��V��QG�Ѐ���!�٠H��j�UŃ4H8ꘐ�p3$�U�䨐�X��MW��lZ+�h:�r������x_˸`��^`�*�q>����ue)��?���S�I�D($Z��1�� �U�Wb;/�:K�!sv
��V�k�Y��C� ,��U���h�/��!M"�Ŵg�|!#�?�Sd�1�f�}:�B9����%<E=cT���f��՗���N>B��$4}�AzidP�Iu7���e�X�!fػ��m����v���	Y܊�W�4:&�z"dV`�#�6M���5�Ҽ���G���Tݭ}��~b�M��^n��C7k�D��/B���*������J B���@D�h]�c�.��E+�D�P���K7��>�n���w�L�4
�$=n].�ޗ��!��	���&pj7ןϝ�t�BC�#؎�Z{l�f!6�/�3 $
2�b2MC�4;^t`�*��b�ɗ��Hu(�;Ґ�'�{��}%U@��9���O�!7'��JM���.u���waI� U�()t�BDۏ�-D���U'.��|�܃TYU$
p�V�RG��x���T�䥫,K̒�JP��i��>a��F>9w���8/�u���(�Z`�k9��[+��!��J5�k>!��C�����b�X� ����kb�b�1�HS�[�����D���V2�y!(���l���W����:u���,w�
���6zTjY/*�6�䢂$R���oޙ����t�c����AtG������G���9�_��_ϱ�0�a,��L����O8dKq�.����#�1ߩ�Ę�P�occy�Z���,A�F3Q���2��<tE��p�\�Xg�1DW�2���A���w��yjX�HU��:E={x�ޮ�y�8�����(,�f���M�.	�]=ʅe\��)2	�oh=�6�����h�څ�3JW@&Hy��E�¼�1ʳG��L�����!�L�M~����'��hK�_s Ua�F�:~= a�V����
K/\�`^  �����Q�"1����tgt�wy�� ��w�!�90����A,P��N�s��U�'σ���k���:I@"�+��X�$_�=�%gl�R�|S{�x���&.�yTv���J[|Em�v��g���2���~Ȟ�y���$��a���1���wC+�NϷ�g�"i���"�j�6��Y=_������Cqd���FK��S���S���HN�Yn�^g�*�V�@O42������{A���-�$��a�ܛ��VF��
���⻱���!��SL���N)x��%#��c
�|�A4�sB�.�V��{h�5�2��`V��i��K$3�r彣 =O��9�4�/���������7Ê-�� �w1!m��U�'�_��Zy'��NY�ܲ���)�F>x]��	&��A�Xkvx┱1c?�؈	��G�It�h�g���h�x�Ij�W���
">j^63 �k��D�7��*��m�A�_���ʨDa]��?��}��wROf����7[���=aj[�)	2��NC(ɫɑ���l`���eS Gi2����o-!}�-�tU/��H�@nG/z!뺯���5�&,������� �c8��4�'ӿ� ��TwQ�߬�T	B�8�u^��ٚ`��0���0�}�*�3�ԩf��<�h�oǁ�T0 ����n��X��	��C�&��Z�m���n�U�~n���p6'�j�cv���Z�/��s�-�v��H���I�rl��� N(��G��Q,׸��ϧO��Y^1��)F��+np�i*���#z�O��5�h��{K@���!�}ċ7�df������6�����g�Vf��V�6��.�z�	g��__�.�ߴYȽR2���SY�M �����?b\@YQ+~Q����ۗQ������'>Ir^b�9��Ah!��6�hN�^ً�®��ͻ]w?=I8���i��V���$�+�S�����l�Ĩ&�[�w�l�����C�^���M��*��K2���������M&����ݬ>�Ԍ�^�?u���',d�[�ru}�Σ5�h9�O���K������\�B+^���W� ��C킂�
�<��g%*,�%�?���|����q���S�0xq��ޓ��A_$���|z|J�h������-����p��K����SK��K�P#0����Sr�Ր� H1�P��@+fN��K�
,��-yL�ZU1J9}�����j���'5������/>����B#/�2��] ��?Ǐ�^5wn�C��(����`y�Pn�$��ڡ��a������C�4-��@�5B�^U텾$Мm�ƪ.&���Sm�z���F�O���z|�,�2b-�;W��%���z�)����1�U'�[��yǍS���=6�!A��%����]����.Ke�E�h㐳����!�A��S���/�/j��Ӂb_ g�'|��h�D2^r|PM�b����p��<r}QV���L��h��랛sȕa\������]�Drd�ρo���<n�Ho_d���FX�6[^��P&g-�����ߓ��\�3L��1O���|�2��;1��;�I�
��
��k@�t ��mprzc-[��Eqg�'/�8=��w�Poy�7�J5�ɂ�4F�YT���>G;��;i���]��`LPZ���u�V����\��P/H9w8�XՊ;���e���� ^?�s&��AW,���,�cj�98��&�p�ח�7��]:gȼ�9QW	�8�y����F.%�Ƈe�A��y1�Ҹ�N�Ԯ�"U:I���t	�/6�@��N�l��#㘥�\w�g�KJ��)!��]�'�f�J�:1�Z��� ���6�rj/��~.I7aUٖJ�7�M�AW$�J|:nͫ�W�S���"��l)*h�A]9(��㻌� ���X�Yӈ�+��1ac����Ǣ��\��h�ٵ��_<(��bM�n���+q��(��=���QO����&�>�������\�xW�1�k��õ����5���E��W�Y4;��� ��w�x�k����zߵ/��>�ؾ�<�L�B��5()�<�����禫9��z�H�/ ~YH.I�~��<�`���ӡ��"o��;h���O�ݖ:�j��l�X����'O�{ɾR	��6\{�aT���[�_����m>�ym�����G�@����!�Z�ѽ��{ﬧ��_qb�[�@��8��PCU���O�g�>4)�rځۓ=`,���vͶzw���P��O���G[��`6�[���%[��&JֆZ7�Γ���.�C��t��۫�B���.��$��%GW�C�A�_fx��BYj`�f���BMt�� ��o[�F������잺T�o�+�@pB���������9NMX������wV.��c��ﲊ�t��(���7l-�ɋ���۝�QR���D���*Y��8\<1�z�|r�J=�8�I�2�9�!��C;��um��>�.lw��6B|�>z=�ܣ�Uآ�����o�(�Y���v�8��bm�}	��\mXdF�ʛy5�y耜��\��Ý�V�
o1����^tj�YE�/��њ�JR!�h�Z���!Y�sq����d-�wv^���4��*��%��=�S��R�=���N�B��Qu��B���@�(/�� ��c0�7{��K:P�.�C1���0�D�d]�����w/���һ R��!�*�BS�uOV_�n���
s���O��f��8[eNey5���	��^$��]��cNP�z�Ⳙ��s_��	��6#�/|�QY6��(�ضЎ��3�RO�c���Ю��?;$G!ar4�v��A��3�Ҷ:O%Gw�mw�C� d�{Q��ƕ$�}lmO뾾ذ�h�$���/k;�@�������Ĺc{��� �t�h[���[�gy�h���`K�Em��΄�g+5߽ど@V�~��?���*.���%�.:F	��r^)�f�-j��=�7߼����
�!�@P	�/v�эc��:Հ,GU_�x7<��(
�v�]�!'v�)��3��>�b"5�v���G�21�����I�b$2�E��>�t҄
�3�T2��դ.�~ᥙ��~�%~G}�F?��8��8�$��ç�:�+ݤ�ăHj'��Yt�&B&�������%K�%
!^_4��ʇ�[��ȱ1�M>�v�pr����S_S�n5���G��YË6�m�a�k�rJ�Zǆ��%qcN�I��9��2��Ш��[X�Zl�Z��N�i>/QV��T��W�����5DE����kd!n����E�*�@"�qA�a���X9��D<We��)�O2M�x-� �#�>�p��#u�eT:dx���,��Z�y�v�)R��Ydi��%ldH�ٴ�%��M~� ��ʉG��V��c늩~~���۸�E~q�?��,
_��V���0U��Ӥy.X����+��-�$R ��D��L�V�e���>I �ܝQ��Z���� �5�uJ`	U�����PR+�↽���T���R�T%�[�~���a�6Wl�]�����U�����.$��y(�t�2�@����!�^@����7x�?@���^���~SvO<o�dK�T������@H>Ѩ�f7��b�EC�د�l����ze͝����-o��:���ѡ�Pú�րu��m_�P�e�� B�����Nh�H�mz�'ϻ�q�{Rl��Lx�b���fk��$6�7L��,G�����{d:�Y��]�1�h>�]Kדx�uY&�!��>���=h�m-A@x+E;$�s��F���E*��]=I�wp�p��PVWN�b�s���'y��<�`D[pUd��^3ICo�K���7:����"a8���Ω�t�c#Ne��[�LG6�J1�#�t��j�L�r��m@;�[Q�2���&��P�a�p���<o2$���_�I�'��%H����$���G*�t)�-�4_���~m���f�L�l�F�"�5�/)�e`�"4�;�p|��Uß77���i�A��<p�����K�vv� �ʒ�d��l��!e��z��*e^`�$vk4e�ã�)r��2����Z`9M�N	n>u�\��`�p2g���oχ ���T�#E����zWv%s'��nv��R��=l�K6E����UA����z�ϩe�~�K��i(-�֮�r������H����U�Dl��8�V8w�
n:�I9��7�P���7�,R��Y���Q5������l4Q���b�J��7R��Ү��Z���ӊ�G�9��f�;�u��{{a���h"AS�Y�����z*ɍy9�_+�d ��ڭgW������(��՟��x�Y�t84k
�s������n�!.�#����_>�>#��qTt$��vP�#����k���7���r3t?]��>z?ԭ4cI��X�H�3�\Y�_�#�ػ:�L�?�77O���̟e�Q�}��1u�N���R����7W��t��������LG(�0���*�d��g��l���;�	�F�IC�`��l����� �Šaw2�ݜUߵ0�4�ډWo����d����O暧�ɽkU�B&�t|=7�E����xI?ƥ�
$��·}lg�~�K�_8b�ߨ�ȯ�����!��J��w�6ڂ]2���k�ee��wݘ�[F�|��/�KS���G��^�d�"���{��H�ʇt����:�v��n�Ꟛ��T���T �+�E��,�[�9����^�B���7�����x�h{1Dz�O4k�xn�S��8���?FDr��͒�&��X����)�@�A�̢�x�	����7�Ͻ�B���ps �̯�)׈A;�!������3��#����mi4����G��E��~$�F�T��.�wU؉FP��t�U6VQ7��!���y����C,^`��2Sv�Yu�_σ;Eo�<1�\m�b�]��"^$gs�����N}v�߉��&R1�oFQX�)�4��������eNƯ8+=[�;�)}�{��*�̈��'���6��,dL�n�DI0���轫�|fLr�ǯ�����G �ʼė����ⵀ���r��:���l�$=�d%�v1��U/� ���2�oKL��iW*hp|1���A�o'̲�h��~�캶G�3V@�2��ι٠˱�K���j �w0���j�v��i9D��ɑ�;y�g<�)ݖ@�������Q�����jL����!f��=�;&A�G�80�m �����ڼ�Iv��s���'���?�����{y�9�>㌻)B�QPz�1�	��34�=��&�݃���
���`m	�8;�<*Z�_��n빊�tT�j��xh�E����5���ǧ-���G�k���%�y~I�	+���X���[|��`s.+?ݶ�(r��n�cѶ�E�����s�L5��]�X.텟��A��%��d���c��n���[m/^y�r�^�[ιi�2�6��\3}<�_nҺ�'U�LS{�=`��4$�r�ɺ8�p���i"�/(�&ƅ��ڱV���p���-g�	;f�cʾ�UU���2	���
so[��ٶ�k�O�2��J|�����"�E��~{��k��P�����M���HB�s�����1~9{�@�����jT�w9ͦ@Oպ�~�:�liJ����N��T]��NoC��?O�{ec�XG/���8a��59�PnN���c�(�y� �)��1���@��2jV���ǉp�[M}�~�֍���z��sb�?Gĕ\�f�I��*O6��&���LY�x��M��z�����-E��%t:�4]�z0��c`������b����/z�[�U���'v�{X��T;�6i(��`|#�%��f��aG��I��Y& 7g����U��ӻW�V$�-|c��s_��|����%8�#�o2Q��,̯�z��k.���|��>p��#</�P�6�~�"��ɐ��̨]γ�4IWI:l�^�q�m�z���R��q�!鰄�3�?�����,�z���82��#�rB	��D<�k;�`L�H�}1�����މ]w�ਜ���;	���Kn���X���l��d�lag�b躃�{o�N!h$�C�ˤ#�?�Hf\m�Vs��	X�������u�g�:����F��qM�%�.)uK%�"��4@�@9�h��0qW���i��`��Ki�8h'�a��E�f��iܱr�}�{���~�!bh/��n��kYg.����}���kw�kX��"U��	|�JnǸb�� I���I׿K��WJ���P"�F�y��ԑ�Y����<r"f�bg�78��8�3���`����hI3�q�fY�OZC���8!@um�w� ��Y��%��/l$�v�PS�n���p��W���P1AH��Σ�3�(ݫ�"��Ƞ����uCP�x���E���@�����O�F;��&�HٲrH�"���O<�^[�̸R�)[3Mx(���'�v��������:�(h<YE@E�����t3��쌮�!��&�K�,zz���N��Z�#�gmk�y>�0X�k�h��e7�G��Nr�`�K��?DH��a���͉��΃�zd�*b�r�/m��|wvI�J
ޔ�x8�hx*J��7��6Q�Y	F�,JZG{��1��L~dd��(ei%���� �8�ZZ�p�츸?�5�?�'�7I���(ZB#[,RtÎ��T	kA.ac���z5��xr�T�����鮳Q�pAV�E�ipY�]6O�C\�M���0��խu�~���!�K|2�믁���C�e�,$��M�?�=A���K��)����A@�-eY���Oi�{���K����d�v�ѝ��[��~�v�6~�x��d���߇�U,.An��^��;��(��C��υ	^��t2�j�$I*9""�Y�����5]������
?���@�IƬX�=v0��Ũ���0(��#X�Ҹ�����T��^a�jQ�(�7_�{n��-����_UZp�:��E`��O����h,L�`q���'q�9e^hUj���?h��"���rCHo��@�e�x4�2 ��F���Q�*�NLށ���}��z"���T��-����f�� �<�S�W��@���x�oZb�܋� {Qd�B�%B!�-�����,� ֌[+�����b�K����H���nbۇ�ѓK���D-�.�����ȫ�|C��zs��Z��xwtx� ���O�M:B�� ���{U�/<e�D$�3�$	�����&nR����]�H/�h��������N����R��G�2d��¢\�c��jHC%����n�v#z��.�:Ƶ���ם��X��d W�҇	z-�9Y��1.j��4���{҇]�!&QT�&�u'��yf��k�](!K�܍���� ���=N�M����[�`\�WY;��g��>d��ﺯ�ůsn�B�ĕ&�iun%Dʸ噅R�U�iGÆ�\�Z)�ߞ9�R9K����5���tw�`���M��O��Q����g�sNst�~3=�Ϋv�M��[���?���Ih�+�����PJX�Y�n�#K��fXv��15lY�T.��?#+�v�h��K����*i�� v��k�M{+�Jk,�9,RVR ��-%���)���{�d�0�-l�
�ۃ1_9<b�W��v��R�϶��Rd��S��B���R$Pfr�8f��<Ӭ�����C��7M�1(�XwJ��1%y����th���u�����X��Y?R�2m���ô�؝UV|Pw�g;��o�� YvH�qa$]B��-U�����1����LR�ET���X�҅  �rH/�����؞���SP�HmC���Ɓ�[=V�cm�	B���'wJF����YpG����?�X�4G���px������Q���G6��W���ep��6�{�J��P8��RxbQ{���bh�V0ԅ����/���-Aw]��ǅ��Sd�kv�����2��m�
��Q���YW>t�%�UĊZZ�,�Wo�g'r+���2���A���e+�{S�u����ސ��A��Gr-W��ϗ��H���S.�Ԗ�:�x>J�G`d��*�[ŅK���h�We�=����@��߄� ��]�F�Z?��"NUVˑ��CKxP��x�8}%M��b�%o�LG5u�z��w��"�;d���U�z6T�Q7�������<���AT�W�%�;w�X:i�c���M3���j�1X�Ў^ȇ�����q��'ruסnU��e����L����vx�	�������(�^C����->Թ���lW~�?�ݮ*�i��39��Z�,w���.y��l5 ⽇ �w�-pa����]ttvy�K�x�&��sU����6�.ηx!Lo��DU�������Wq������
�،���*D�Q�)Ҏi+s$%ԡ�>�}*J%<!g����)� ��uP�?X��O����-��<�!'=AuW;��<�Q*�8ޟ}�yD�K�؈��uY`.ZیauhKTk���*�V��Bx��F|���Sƒ�Y�i8ΩT�6p^��JRڵ�9�V��5�*[����{�7mnbz�}/K3��	>v�CL��3x�§v�sבs��hĠRd�H����n��p�.�_�*�޼��)Myy�|�����H#&U�[҇&|���!���+{���t�~��#$]��8)P�I��]�^D�s��~K֖�O�jM�߶�OM�)�XF�Bd	�Y)�PX�gÆ���6���+�k�=���������h�E�yj4�sz%F����D��5�.r���\��d���ʬ�q�r�ڢ�kO2`������o'/�a����;v����K�������/� ��P��י��y�F3to�uU�A/5!����EA�7�ڞF��n��pH̚�0u�:�g���tR%t�����˥�!b
�ޏ##3��uFe�)	�ݕPt�J�/�ip���Ƣjxת��� %Z�-�7k�x;gh� :�� �P�+�"���m,�n|�p�=r��#�a�e�� (
vS=�W����l�K���0�Q%����H�6Hk˞]��Ѭ��Ʒ��ɸݖ�2��%F���y���9|�L���O}����Wƥ!4bQ@��l��Z�ڞ��fq"���u4;fK�ti��6gH^A�hq���aHN�E��ݩuDM�%��=I��x��mn�Y�*���p%��3ȶw��C�6��H�/&Õ�*�	v�\�23��j��%��9��p�����]E�(�u�ݎE#GJ�R��o��xg
k�-пw�����@E�2d;͒~D���iJJ_��ftȔj����3ɘU|��V1��$��UnHk*���Y����O��яo��(��O���m(���\#�[ �3�&5�P�Ν�x�f����T����S|;׌y0i���
��pƨ����_[#���ovS�/�ʤ_/ϰ01�=5DÁ* � v�D�]o��?9��
Ȼc��Wj�TtIxֹ�D�)^������v��:�g�=����z���`6&5�=x*�����G<� /_��V,�	�� �㽬���\<[޽�����C|QrSw7N-�\�#�+G�=+��ؒ��z�ŇI��&�.b����8�j�����լ(W�+T��-N�����'i`^��zMPܨ�Wa�}���_����e[�����"p.�dC����~e�iݝ~�=7���fSp}M�\�n��wﾄ$B�؆�jVgۖי����_�og��'�n�I�Eޤ҇K�3s2�1�������(τ~NI��m�mj݉t�E6s�	�ð1�!��6��}��D����g�b�����l��R�i��6�e�\14�o#.)�	#��]j����E1�)ÀK���ɚ5�MaRk�Wm:r�@*�2��rUB�U�-��u�w'��U\���ǿ⍿� ��+;5Og{6\?�k�V/�.�z�<��r�B^l3.��A�}\3�e>���"����S�x�)E�Sf��Z~
��2g��I�������
�͔�Mg�'��"�O�|_��_�%���{���ԏ]��u�{��VZ�_��g45lV��w���<U�[���ΏM�F�]N��*�ޢv�ؘc�{�� ����^C=)�e��7G�_���;�8�|UQN�w�7s�5��g&�v�%��v��|Q�a$�X��I=���[hlu+/�/�91L���T�m����n�"��'�}��D3@�]y'o�QΓ8��Ǳ`�y�Y%��z?� ��0zJ�>E<������\��8�"V$2���+S$a���ޝ��WZ�HUh�^��G�ԛJP�w/�����r��/�+)���v���$O��^v)&��nf��&9�RE�����N
f�S��|������=��k
���]��
��rR���N���I�>p{m�!�"Ѳ	`&��*t@܎�wZT�s�ZV�3P���P$��+,Ɣ�t��`�ZS/��_uS���-σ��.C�M���7�%Q%�=�㊘F �y�I�S����W�
q�8"�0A	h鏁�M���~	��ǟ&j8����{���AT� >��D� �N�>�p{Q?��*@~UcR$mʅ��P#�enC��P�!�Fх3H{ C*��oq��g&�����Ɇ:�B���0b�o���o�ê�+��^a���ǽ�p�1k�iJ��Ƿd�7LM�JҨ���=�D��a���H���Dձv�B�QD�=��a��&;� �{KPJd�6gzD�җ�!���{���D���G�>�ݓV�k�$��h�y��V��ɵ]�ɱ��GKaV^{=@[��g<<�W�Z���5(�P�5i��gKIj�l��t�/@�n����)+�E��EB+�� ��V�e�+��5q}�Rl$G�V\��\�IN¶�����L~�Mig��6��M.w<��l$4bgj��ǟ���"�	_��v�[����%���xȔ��	���	�[�k�8:���.-��j�0*��"����(�Y�~�>HW#羻C:mºŋ�+>��_5`��ټ�U��Q�3!���{v�Q賹�큥6P����&zMެQ�{�ٜ�Y���o&0b���f�FZ��Q=���Z07���o�}~��G�� |�!� 2��T+���R����6]��5q����;\-�*G	p-g��'eC�s�iQ����37�o؏[z��ksq\"m~���m����h
���d���G�>L�x&9V���3� �!���^��P��)+D�����#Mw�~�e=��҂h59t�Ȟ��o��Ef�Anx��:9D�ax�Ӕ�15=�}��Rn���b_�����+�5�.u�2߭���o�9U���)�s�8v�0Xhxv&��e�ltO����L��~���:�<��`C��Q����$ύ�����K��D�Y� ��wy�MQl��#��7�Z˥�`�4�ev��À8����D+�e�,���-���9�ab�a��O�?���a�������VD!!��?�����ڥhGg���Q��)�k�@�ۯ��c�܀W�"6n_�х-�#�l�0��5��c���������'o��xj�E�x�H
�v�i!����H����w0������(�?a#y�j���eN�4s�8�~!.e9�V�Yr&n�g�=���]���>�>�·G�[
�wf�1���h�u�e��=�J��L��I������� bD�ʸx��~ �,dv��s�k�qI �S:>�	���Yy�FL�[
�4.���ut>4sΤc>QM!���L��`]�2Ԗ�~^M#�Q�`��١��)*/C��:�x�z�mj��l�!�I؝kC+pI����s��=�NGw�1�s��'�w0O7�!�k; �F��]��o:ׁ�����+��K���ΙlÇȅۑ��f3�ay��w"����k�����Ֆx�O�mKL[N��� �Q�s��&O(�/o9��ѣ46�N6:p��#ء��k�DW>dP~T+"���`�������fMk���+,�<kx�7ixGU��	,�Mc��S�{|��w�
��k���Lw\���� �,�RQ�.f�$��x~���6�}@���Ҍ�u�iH����Խ=�#z�_I��a:�b��h���Յ�C���ग़�^y[4s���%ؒ�9%�XG@���H�C�;�W��I?#���;�@1Ҝ�d�?F�N?L/*�#q��C��nx5�I��r!0�!H�� {Q�#+�u�V���?�Ah����l�V�.;Q>�
�����H���;a�3^�3�bTAe��]
����%�u,�o�U�I�T�YFr@�y����J�
�����G~kM`GU'�ق��F�P���퉏p��$��@/J��je��ѻ���f�;��F@=;5>���򪧿���[a�>�Չ�,�p���s�8��C5xLI�7�fo��(I� ���W��~��;�3�ea�\붳i�n>����c���U}��D�r��{�UC�8��<�+��d-���$'>��_�p�͆�jQ;��(׉=D,�xE8t-@�7���e��r�O��U�Y�m���@��LP�.	����� �.�Wo�y7s�˭�������#��O�}���w8N�ڵ^��@� �w���Ə{8|z�Vջn��u�Ad�\$�
�jrD·�,OU�&l�̶��'i=�zx��R ��1}������:���d�B��:0���Ŗ�:�)�&���1nlK���
��#�c��MMG��>� �l9&������C_���Q2A���Z���]P2��̢��#� �v��a_�P���J
�[r�_�Ktl�*سv��Q�t�h��iX9GC�P�` XR�6G,��Ylwq0�����h���馯ڼ=��(pq��l�'��t"ٽ:�wx�S��V9iʏk���u<�e��w��L� 𮧷�d�1Eƛ��L�3������gq�ڊ�֏rdT�0���R��?�j=�)��{>���~��Q8�.�4�ɊH>O��1P��}�Ã�i=09�T������*��b�w��4u����y���l�c']�"q�w<Z��������$S�huF:i�O{O:Aih#�&�x3�A��� �H���
D�M��u�-�k!�|R&��ox'�l�&,��mR_�#\$mA�O�6\����[DBsu �*��澇י�HKW��<�҅5[�d�)���۾�����2&8l�wl���-��ƞ�dI[w���B�S�_2ր�Ka�٣1��Hmdk�A�+�_z��"dH���3-�J�@ɛ�r�����o�S`�e�?\���'.u��=�fA�ǥ1���V[#A,������j$磌��C��W4\B�.�I	N��c�|o�[���+�KNsM�O���i&�񟳣��ƹ!�NԀ�ȹs�h��U;bd���^kD�����R��]{;vƅfd�-ʝ�e�������-�b�[.������}�]�1�;XP~��c���-㳊BU�T�ЌP��SZ�Z��}b�0	�D��_\37�|xq.}O�%Q������Co�y�k��_]:(�aD���K=B7�}�����-�@��Y,2
S�~�WGj(i�"P�iz�\O��:�Q���ǈ�4�5A��i�)T�)e�Ƌ[L���]�^U8�-�p����l >t��_G$7C޺���O�ɥ��!�3�U�8�5����|�+�����;73�@�[�]��VZ�5�*;+��`�\m�)�;F���g���Y(������&�#��[m��)ִU�Hd���'�р�����_��uxA�����4������x�ù���̐��d���7���&xzN�Nx��4\�D��H��,����2�.���`E�%�"�F����Ppw[�h�Fg\��f@���m���ݔ6���D�T|��_х�\�t�Uo��֒ЕØ⒑�)De�2Y����~��m#�"Fl��;�(���ϦS~+�k٢����@�8~^����LN7��1��Sw��y3w�kO�2����t�.��@��?�g�6$[��{���j�M��_�� �/D.��P����t�Q>�uV�J(�dW��	��5�����Jk���
3.��l�a|2��p;%oޡ<Y%�b%00���AY��f����aU���{L c9٤���%v>�{vub�c�'h�w��wW
DF�髠1�[�Q��z�2#H��y�ݔ�q`��v�+���<ěL��b�J{�z�#��Ff`�A�f�\=��e]�;��㲬�����to��O+SP՝V�M��u�Q~�ȕ���\�6��^ΆI��?��,�����[~���&l��L�\![l{df�
е���nP�5��\Zm�1�Y���d�3y�_$�����8���׈Ȧa��u����s�9��7EQ�ݧ�/�XX�"RP<ĩ��;�
'--i��[��8�2�ؚ%�z���ә�=�kc��g'�d�D/�J(�1Ү�!tJۚBrݱ��9�H���pS"���*Ía�}�+[0͌�(j���Gw��g��W���v��X�St40*�-q�M��޲z�*ҁJ5����q:\���͵�a�0�H	�_�6t�Kv�гrs�v�)-,���L�|���
�XA�$4�7���?,3�5���A��n�rY�+�s����.e�K	7n��/Z�0��Y�A:�*Wy���+��M�J�q��7��n��K �J�`�*�=րp��T�~�>��:WWE���3�fZ2|Ҍo0N;o������i�%	��o�����G���n�S	�ƿ��.y��r.�~~EM���N�5o����6->��B�T�=�xXU/0�5QH�j.uh<���R���SP�:�|�١sq;�1M��֫F~�?&;��6|2&m�6U��3�8�m���I��
��wEU��[3F��4�l	'��O,�x���;�:�����7k7c��Y0^����>���"�VҾ�u��`����=x�̞�э���{}_�>�o���a��^�W4��$#��!�ì�e��,��"�!�@�TD�:~CN�`��8P���\�~k�H�&�z�(�aZcǫ��gI�8���^1Cl�&"���&��+c�k(8��hI��8-�]�~�{��L�l�]��Ya��X��i�{��d��dQZڵ����}9���rbײ��),<,G�;^^}i�ܼ�9�*_@�t���#M����ϱ��4�M�\�i���W�S�?�L'� ���I��:��O�)܁~�x��"������� CH��a����aY3�Xq�����pv�DFWϸ>���-[J�m��}$Kg�a�K�g�?��5aV&��!��t��I}�	��Z���c���bƌ�lji��V��;��jN��5�Ĭ�r˗T��pօǑm��)�)��sj̶(�3�z�fL"d�����CKF��^�k4F��!�m����]�(�pp�<e"
¿Ʈ��dt���x�ڏf��2a-E����珚
\���jB�nꞌu�y�k�g�.�t�ZL��XZ��Օ����O'F����� T���3�9wd���힏��˝�H��c�0}���P�R��-�~���W}�<�*%Gy���Q�4YFd�ш,I�lW��9Z�i,��)Ȟ<Ş���-��&ּF��;*F����a��i谏�,� 	�i��m��"�m�����v�z���/@ҍT����T���5Z;���0�\�\�b`{���㉚b(9UI�R�����;Y"�U������W�*��ϭ<�+��C2��_A_�Pc��P$x�U�	c�`�Üz�"�9��u��*���Qv7��t�H<u��n�ei4U�g�R�f�N�����Y:PV�h���G��
`G��j.c���V��X�z7����20)�`��j�m]��"�I��m��Oj��;O��T����q_Z�%�G�U�i48�R��龸�D�����(���m��A��H���Ppp�b�WR��3)�	nru�j;a-8ξ��#�Lc>���Q�\Quy:H}�f���	`��Jt��k�����A���G�6#���;��Ѥ��B��.Ʉf�ܗ�z�^ͱFM������J�	�>�1.;���۞+�c���G(
m��?v�Ng[^'*qÃS%vB�_�F��Ww��jy��.^]��������6]2�ی� ˳}M�dɡK��U��"Ok���TU�G�b*�@
<�9��(� >t���p��O)}�a�#}�ۆ`�Vj$���$�o$�}��V�}fNQUN�I�Wi���P������.w���ܭ��1���9��ؗm�~�3�2�J��C#$��p&��&D+�zHl!)98aL��|��v㈦�SqD\S8��k�/���ڲ!d`��c�A�԰�_��V�22vu���ȧ4�r��(`_�:�&��]��;W��? �N��J��|c������I8�&��k<��V��t�C8�s�/��	twX 0�է����At*ѓ�W�T04@�W���k��w/g�#ر���q~��G�3�%r<H5϶g|ρ��3�L�݅�F����/��e� �v�7L��ۏ݊�ʂf${������%��%�~\�a��&����!G���] �������}�1ݬ�9�)�N� �t�W^ T���V�!@�=���d:�6�Z���������Y?X낅�]x:\�ٿ�:���m �1��v� [>b�MZX��;�l9<����ھ@G�C��\�@�Z�it� ܵG�v���}�!YMM{+ ��
��A+��0��R��m�kė�g#s�L�.F�%%��g�Ě��&��`���
4-�-G.zq����Rj>c�)���0����*������D��eI0���k�Evu��^��PR5�P����e�D����G�",�Cτ��:o����C0�=�o�k�<�OP04�.��t�,�������%
���֗�������&;�@ed��xB�UY���8�ub�ŉ�B�v��w2�»8�gn�Ŭb�c5����2��ڝ�����`,NukUv+%7Ib����n]~pe��з����!G�Q��'RCB�Pq���m�ʁ{�M=y�n�)��3�oDf�G ��F�������ʁ��i��4�{�;�r�IG���S&;i�6�~D�m�g@�� !fF�|P9/t`��1�������P����Eߧ(��_��+'�^��L���t���(��N�#MJ��y����^���>�&PgV�)_���ZL~W,ѐ��M��nkٿI�D.��E��C�p%�9^�wAg�r�$��3��fm�뫛j��i���L׽G}��j$@��b<��*G�����~	�6y�4��Ǯ8���L�8*n�$�E���ȵ�-�C�Kf�
{�$?�_��1���V�p;g�aV�ȦP�ɼ_+J��G*6�.��K�B�i#L�!}Mk;�����e�j��he!SP���H�����ncǄ�R>J��������?qp��]4�]tO���G9����t��	��j�[zl/ߖA��[�>ӡ��F�G����6�Z��'��ͦ=��x��a3m�?*�e�O��~M,����f�Y&�UvOC8��}o��wV���?�m�wmFf*⮩����ٍ���T�S���{�D&�1��h�kq�`��]R�WxP�� �X��ؾȠg]�{v5�����B���M�6���T`'�N�3;��I�W���6t�sS*־��#��`��r)�w����6Gyd�S �� ��1#uf�1�1K�Gu�\��-�g��;��X$�=���4|�0�^V��M�Dvx�R.6�ч<yY\��6��
�*?^�_A�� ��&.'�K+���l�����3�T�����+���LѿK����	�@���r���NX��X��yt~	��4�'b�0aT�d��`��~���I$���̤D�T*qW>�O?�*�}D >a)c�p*�H���D���e��(�*����p�cI�B�{�_vB�%b'�rL�9��@���;�瑁��%-jWn���(1S*�D��9j��i��_��Or��f�+��ez�x��f��tpQ�Z�c�&='�Kx"'gi���� ���[)ԍO`�+��2?�N�4zR��n�7���At�.�E�;`��Zk�[�OD�WKjZie~ET�m�P[MI.F�~4��<0�cz�r��=6���/&sPt�a �%�f�Y�4�E֩8b��+��d�q�zC������<�vZ�X�X�d�����Is�����~�ܝG���b���+�~%�_��>��Zh�J�W����T�b~d����oO軸���"�8#�ӋW=�,Y���n�	=���DA��:a���+�b]���M���Y�T��<���{�"<g�$C)����y.��#���weXv�ޒB.���tj�s�n�:H��v«H��>�f�)!RU/6��a�9��7�'�3_��Qr~�	+u�C/���W�[�D����i��1Eg��*�my��i6���̢��g`T������Z��U(9�,��Fַ�%��]'�o�R��n0�����.5�aȟ)�jR?��xkv�O-.
�\����封�K�	'�D��.���tb50߬ȶ��s�Y��R�<��!�Ѥ��bަ��\L(kto�(k���,R��ػi<���}>������p�1���$�?��U��tQ)��9��c��� ��x8P:����ca�t�P�)7E"��Qi�;o��|�)�|LmrYc��]�����g�l������N�~ʦ's�lp4��Bt�ݜsH���3=i`;������ĉ�M��Wf���,������B%1̀�?�O��@m�/��,��#�z+Gt���Ȩ9O�*I�b��Q$~��%'~�\?8LLgT��\P����b���|�P���O9�����K�4%�9�|/����2B<�uB���	�E�	�F��G����h�{�Lξ$�fvX��?T����i�
}P<��p�P�����9*�qC�ɲ&ą�ćU۳ܡ�'�,��U�)�fkgZ�T�����!}��G@��ӦT%�ZvWo�0d˃kzHu���#���3>1��b<�pK�ki���^iOMM|�������OU�ж��0�l�h��E��t��q2��IP��ڛi�s{����/d5;$߽͆G=��|�
1g���yM)_�	p�}�n���De]#-��������o�u2	������	�i5�d��(B�B�}�7�A�"�<�3��m���/���&�0GR���*=խn�ժ$Dt��,�+�bg��N��$�HY�U�h&E�8o����{�6)M?���^ހ)���&��<��L���x�����������L`�]:�L��9-���'�u}W��;;�뗵6O2EX�Í��S�+��"�z	1�B�CL� 6>Rl�4��99���{(���0	PE��<h�����f\�^LN�^E!>q#(�6ぜ��BZ�+��d�)D�x4��钇_�'�o��~��Ź�4�-�v�j+Ьv�Y}l�k��kɎ�K*`�k�z���=�}]��q!�끅����-�S���Y��~��<s������|'��
��ȞTx؂������/d�gBb� Y��=�ˁ./�O[����\����e����B���G�Ne`����s�+�0o.~5vRX��A��$)�~����ҩ�Z����J߱+�>t�G���<��i��]�Ne����+�e�@Lئ�����$��A�!����.3wn�N>ϩR=�<�!y��)��4G��bm�M��j��K�}�}��#���=%�2�m��DG�,�ݒ,�vwq����,����������������sy�?ct��T��0L�T�`y���벊�� �#�Ǹ�u�	��5��ױ3�ȏ��܋�Y��f��hƱ������a�ne;�h-�<r��Q���@�1t���d� ��]Y�)��$����`Мs�*�����-�e��t��L���L���r���Z� ����C�&��U�P�TA>?��8�4Wh�'4�r���;z�d�)�c�W�S�y*��g0R���jn�
�xd$L9�C�H<~H���<���i�V��V��5b:Zw��� ���U+v��I�%g���ȥR��˨P&��o��<�P�����󗚽ג���e��1��kk�)v�m�Wb��y�^:�#9�(�k�����tѝ�%�(;�6��c-�k/��z)׼����-����a���<����t��gC\�E�>��b��E����xDh�_vEkF�(�~R�?ֆ�V��n� ݩ�S�L<��C[[F��X��h_A�k"��PA��{;��Ӂ��(l�|�5u#��gw3��r�u��1%;�B	[ʝMX1�����|θ�O�O.�O�*�w���q�����2��4v�<ɲĳp+�V�x�2�y' ��
�d�9n)s�=~�q����X',�sGv3ǐ>`��Ѵ-��ܝn���VX�5��"��A �Q�Ͼ�����M��K���ѤQ�C����Q�2՗�A��~�Ȁ��@��op1WO�D�6��:�-���y��CC��I&�Y�����ǉt'������}��j��c�%zO��~��2"�H.��H�6���%�ؔ2g���L�Ôm0w����/�pv�rĬS���˟�A��Gp��e_X��������1�.b
���3���:-�^#r �`�k!t�пmY�/�b+.qIG/3Z�9��`:���X
�����K�h�$}������P�I�MNad�kf�(Q�P}�F�v�I���y�M �z#a��?�a�A��P�xtJ�y�2~�I˶����!�R?_����1cd�evVY��x�O���,[�hS2=0��Do��Iu1ib��[�>���s�[��/ҹ�WNnAr�H��0��n
�i����"M�B��4�Uݢ􎨾,�7`�-���������ّ�?����vj���+�}驰�3IL|N����6s;%ŸZ6ET�Ən�B�x?�%���`���B�ʶ����6�;�ԃ��l���	��L6�}�u��U��]�>�5Ga���jҋ+.)�A\ǰGWA�HmNx���K�]�;�")�^��p�B�%��zAs��m�q��&2�_<.8-�_���=���j�*��C"�D09'z�.��,"��Kx������^v6Z�YYj��K��`̷�*���xV�:ܖ\
-7��k{ќ]s�m������c�NF�+gr��1C��'b�9<�n�}���o{+�K�P�k��gX�J��G�}]�����cf3����R�h<���c���n��������Jt��t�h���((�u�a���5@Sx	�NJI8��|H���	,�҅��Ey$`�o��P�A���o��#2�9ha�9ڐ׏��"�����4u�oa���̿�&����Wi�JLVHJЈ��$�u�:��,>`8*q������_0�
c��C�s��`4���қ{`B��⼂�E� �\tT�6q�?a4������(�Pߑ꘥VL�j ��]��|�y9Z�X�iyXUc59C�%�oȇ����w,�J�dА�(��^C� �s�M���,}!�!���e�Z92u�$�Әjb�x��sDI�W����>�ĺ�S��գWr��(
���4�u�9�3w26�o��;2Z
>/���|�z�g'Z,|��.�䈉p�x@���F��9��=p:�����E���j`a�?<����O�215�Y���A�j��/ՙ9T=TɧXݵ�Z�Pu�[����m$�Fg��xXn���1��~�N:��q�BݞE�.�	���\���#���g�:�칠{0�[��}g�|��'Ч�R=^�_�K� e�4���!����P2(1���E�ef�p�q�å�BM�[UGO>����u=�Pw?��JوTeY���W9��b���$�&�%Z��uɥ��Kk����\�h_����l���̻	S��d��Y�-n|�~т^HWl���bv���Ν#��j;Y�}��J�`!E4�5�_Ұ�5���W!��eW�Vo����B��n=\Sӄ��>RU� �Hl���;�M�)*�� >yĜ/�fitۅơg�7���� �b�[z0h�?�oM���ȷ��Q0Wr�F4��>�o,���*1�Qr��fl��c}���f��D�~�F	.s�����[7"����lO����*����tj-+͑�\��0	����)!��p�QK�׶Pj�^�(PT���:^+��,�jP��~�fC��x����?�x�~��,,����q���a��@�I�A LD���[;�6��
�u�f$�m��r�㛢Ft�<���*����<ǎ)+K���8���{ʤ�i!g�� ��N�)�-~_O�Х�6(9ʲg������|2*�f�4�d/���86�d$��I����e�Ù�f4�s��^��E2����<�D�Kզ(�O�����Rt)���}���2n��R#c��-�t�Ά��c������>���[]`6p^)���/��r2�+Q����Ð"�L����Q,j&����8���E��%�l?���V<�8��R�Mڒc|�]�';��g~��&]�8�ݵ�ϦL����y��-W�i^aR}tHFO�N�!¬����")���	8fd�����t]���Qd�����q��Ě"?�FE��b�uDf���F~�Π���b�>-��*tc[J�N5�:g��6�ޯl���u��lе�6v=� d��!��v,Ö�3緇�k�4(���ޒ�����zV+�dFbҍC!���������R81�@��A�}7�â�H��:�jW%	�h\@�DMS*$��}���V5P�*��˼�C��sc�ϔS��tQw��E/:��HU4�&y����r��K��?`��g>=�/�E���h�C�O�9?`T�jx�p�=!����E���S������8��q�ݏ���	a�NCB��O�yw3�2@IA�e�9~��q縛�/=�����w�a�����X�B"�ӯ���8`�sLC��m��-d��>R�U��X���G���Ǹ�LxY�ڛ�\�]�-8J�2�A�8�J��!�pn܎w:Y�B��&xUp��q"@�*	c�w�ߨ�^�0��>�����T�櫘\��y׍�P��9�t�w�bJ�#8�H:ۇ�	��|��J%�/��{��%'�����M�M���yѣ��Y<�P�ܟ궉��� 	�p���8I���Bk�,4���YY,.z[B�@����Lo�ҍ�m��A	K��p���/݇��������嬋������KZ�����;1���a۱��� ��|ՏE�T���Ok��6�i���KY�}ML>����ܟ�c ?4C����sYD��Oӈ�F�G�25�fx��b���1��UxOZ���#����3 dZ�Q�?Z�'g��s�|ٗS)��^��W�e��"F�����ܛ��N pG2&���*��]�� �����$�
���~�]�\��SCR	��G��	�������D+�<��ߕL�}��9L�;�t��2~�c�B�U��Eo�.f�Ё����?�ʷz�h�Q�E�ND�]6V}�G���q\���C�����N�7a���xr���35��;]$����b�%�j"�.���fHw�קк-й(�n����'�0�t�Q�ge�N2L�Q���D�)+�R�ǟú�D�1�]/���Ix�{�!�vW��1� ���.�� ��G�o�C�_F��1i�L+��>M��Q,Z�@͓�>���6���#Ջ�rJ�����m_��:�hgo4V u�&��v�Aux�A<� 3��ʸ�{!�<�mw7��S)�#�4`�{���5Iԯr0�Gs�N�'[���@;<�'�Z�����7*�+������l3������y��lz��ᨴ龈�^����`x�L��)E�{`�p���u��*Ծ���?���j�w�<1��e����E�Ѕo[V���u���QaL}�cJYw������A�Y�)��� ��{��H�8�B[���3|��I�ۯ.��+Q�{���E��@�̸���5�v�����Hz���\���C����])��ҕ������9*�vU��'���m��̦%!PS׷�Y)������,[mB;{���N�2FzJ|�fς�´YiG��+�j1�ph�wwĀ]me�sl5��; ,��pW�?A�z3�����+[B<3��\/�<ҏ��O���-�TW�M��E�����<�Z�i�9�v��Kԯz;���)��@�K����o#��+k����{�]&��wա��L���V��X�g�x�M�Mm���J��7�<S��x|����^KW�Sy$��*GRFa�\���Y�%m�r+ct�u�~֭g#5��� ��}��K}#�{t|�}���Q��B�.4��3���C��b�j,��g�dTQ���.Pp�HI�^JNں�X�,���7�ʆ��,A�;k "�}���s]�ƀ|ΦU�It}jµ/:�׊6���_��F[�Ϗ�P��u�g��@	�������}m8�ٷ|�"q�m�'�`��T����l�Bذ�3�U���VS���#^��;W���b�T�}�z�sȠM���<�@���]��#������ʗ�c�e�ąK��4� � ��`�Ok+�G�����8�[�@�Su�t74V�tQ�h��2�!ռW���qd�N���1�} Ϗ��dv$�H���J�a�����P5��.���ٝL#P/���Bipq�݃T�e�w:�k����0`{�|������t*���M]�w����d��Ͻ����	�n�]���`�P�0����f�-8T�U�pgJ��kr瑴1`��I[yޮJ?�3r��\�s:V!� ���BCY�O�-�oZ���c�����X��jJ�N�7�%T�X����dY�y��?��EW椮�^7ah�y�'��f���t���k��'hk��7��|6��
TG�=��lO?bl��$�'�M#�n�e�����,���0x|ݕR��|���I�7�����|�?�^���U[���;)��sa%$��b�:@�T��7�(t�HS�V`� ���,eaz������=k&�%=%�)�v��mE��^���hz�5�-�������ͥ&����^N����FJN�:�;��T��i�鷏N���k��O-:$]ХG)�@�H�%>cVr�u�)b,��h�";V��A��6����@Ի�vdo�ɯE�Y�:�>UP����ZFY����Xޔ��m��'(m�pK8�����R�1(`�N�LĒ��8��B"�R�	����\�ߡ9�>�.&J�Yq�c	����ޥ��#�u���Y;`!�t��Շҗ}Q(������0��q7C��A@G����ki����JC�;&��VxX�[�^7WM�܀�N��Bu�o�I-�Y˄:�E:�w(0zY��� �lu+�lΙ+WV��|f�H ^H<\x6��0(�j/�sDa�"h�&nG���j`s8�R�o*�������o���C���o�
��'���x��{��F�L�H�.	B����\h������E���B5�vr�y2T�iҜ��� L�7T�V��x���I�`L�w˯\5�Ϯ�2�|C�Hx��?��d�M�&��4�n̽���e&8�'U,6�U��R.�A�i���Z-�V�5
�s���M�Te��}�!��q4�Io@
"�M��3�}'��^�T5�S�s�C
�C� R:���eg����&{x«�K�T4���(���/����b�^d1�����F�&`��G�I�ӯ�8)�82� ���sUw>�����E����LX�u�V2@�x
�������+�	������J�¸g�a��tg$��J�;����D����M.���^I7�W�^
�C�{�%(g`��u٤�I����l����j�6>5�K�\l�ۿK��$�>�٠`gPf���yo<�K/�ɜ8�=����޽iXQ��dN9�PH�T�?�L�� 
��;ȀR"�0��Wr8�%8�!�S����f�;H.�Τr9������EB;�p�x��d�1&�\��a_%�X՚�-��,�-Tұ�*.�s]U�̔XRѲ�� B�0��E�A}���P`��)"<���^y��K�0��D=[�w=���!�N@����ۊu!{ ɱ�'h@�,fF��`���l*��q�x-��1� &�nr��bo�CQ´>|G�z�]g�=5 dz��5U=}|���?'��|�[iK� ��	6j��6=[��3�WS���܈k#,$:��p���ɵu���U��h+�@&*ֵ��B'�;h�����GD��W�t2�o�C2�E3W�E�]r�,ϊ~T�SV!�����mKN�R��w��ȴ��s2�29��'wl���u�O@�e~r@���1ANg�Hi�
I���bV�F���35�u)�[�'[*K'�����XI��\�:�E%���.�[|�>w؄��PO��|�[�%#)��ߗDPOv^�V�~��)"(�<
�4�m�+���4�cg�4{t��6�9�����O�'�f2�۞��pO�$���y�W��)q���a�؝n�ԡ�V������;�Ld=��#5UC��霑��?�B`��Z��N��ܻ9?x��I�J�b
m�/�ڧ�ƌ4�j�� :c�#�)���-�X(^k�/]pk����} ��M��q�������::") ��F$Y�o��R�4ӳ�4-<\D�z�¡��InzT_)�r:PNz�O:�(/���ڰ�Jr8r�.���*�A[]4,���:̓��a�3�D�n"+NòҢ��U7&l�A���6�R2,@k�my2s�fַs��S���k�[�lݟi�>@|&�����Jm�i�C����}��ģ}*���S���qS��� �Q*�n���1�����0����r��@�ݑyb����d��D�S��4�@���QR��97����*�U��)e���& �"S���E����m�gH0L2�7���1Ļ��|���Y=u6�.�����%?A.[is����^*�W}M�!���w��3�_���@w>=���O�cؚ�j��>s����ȃK�s���_˟�Qr׀�A�W�����CVi�H�*
�q����s�����Ϸƅ���Y
S��p@�v�˝��}�o=G!���P*aT#���C05A%&��D4�o�/I�M��ॲ������)�*���M�o�7������aT�2�ޔ����5M�Ó��C���{儚���X���5�NC��b�����s�9-Z-�i�����>�V�',�����/�|a�)�4��?g�%f�U�������&/~t"��lY�Ǩ�aHح}d	^���"hv�(�qdL����α�U|Z���������L��nJ�uT�V�/���5�DN�lt��z$d!^"��w����x�B/bp�A=]ݴ v�Nvf���@�
��|Y�)(G�.��l�2);��ah�h'�aw3�t��؇)JɌP3Z�L$C�OTl>d8�w�\���(X��0��Z4���*�w�@��.�I���Hy��+x�(���J�i�Q?)���Vpa�������#�ݱ�6ӌa������Þ�p1Ć��
���	oM� ��s�FF����zDKU|xI��B^��[�$���Zc�p��c�� )�������zhwF.�[E�SW�gy���yPo�:�L��-ܴ$OA���h4�U��!��=�-����_Æ����9�Sib�6��P$p���{�l���4��)��<P�4$����3I����gpr�i�DH����IE�3TBМ:P��A)�؛>w��Y\�O��T\B%m�_i0�~��&��{y�(Z�Ϙ�
~˗�8߷<}M�bb	a���/k�2�^(R�Sσq��eA#�s�XQh��C� P��:r��[�l�s.��:J���~D�e���a�~����ҐO��3)���a���bѭ��*�W4 ���M�S�W+-�É�kn�!̐�䳀��Y|&�Rfb�
���Zj�*��ʳ$�8�ior��[��g��;�T0[�r��աޚlmv��}�6��s��8�����\k�3��٨�X�G��8��� �ڇV�J�a�&���=�oCҜx�{fOy������YM%�?�j�)�:Qk����s���\��Uqm��'�������<��I���F�!&�Z5�O���1j��ъ�D�>D�t��yL�;rH��]b�(���e�b�kO1�d�I�����G����U��[ׁ���H[W�����-��r�3jּ�At	5��5�~�wq�:��3����NM�gb7�퇝��kG��1h��=�Ƃ�Z8���@-�~'�͚)z�����Ȋ8�����i����w�e�Yy�;�/��Aќvʴԋ����=�H��u�Ǐ�L���/��hmV��Y\Pb��g��lf��a�m	�Cm6唥B�
��q�w�*��s�˝���T�����"/�ML������],uu��g�����ƀX���K��]TM�5��CV;3=˫>�n�G�N�}��*�z��o�J�킅]����
��r��b>r�%�f�T
��nd��{�jfp��	9�v��gx(���K�t��n�[I�&�zĥ��T�{����Z��ww�`��U�[�@2���%5]��a
u��	^0��i�cﹾ�d�SԔ39��:�N<I�{m�О�']����)�A�����H<�BU���tˎp�s��+�~ɮ�r�=y�L��"`��"L�H�?a�*&&�ͲC�c��i�	����x��|Q��~&/��7/�:@Q)���o���o#�)X\똒+�h~8�1\^ޘa�q�e��ϼ���z��*o݀D{\E�n��(K-�p�>s}{�w�|�=Ov���X�4]�҂�����r��[9	��������4%vQzO]�-�#���y<�d�|8!ȟBV��qi�f��;\q� �Ao`��ex��e�������#���N<0��	��V� ��P2Y��z�sJ�k	�S~�+��|C���#��򰿙��D�6�b9����d�Z	UՓVã�ʢ�������O�|h�RԺ[9V�?,�{�k`���f���D͗�{�_o'����6b�P�^�I���ʄ�\Sh�՛e��`Qr�i[޲�Z����|E�
�;��N�}�He;�����;	�t>�������M�r�����&��7��M��C�T�X�_��l�Q�פ�^��^�ص�*���dG�&r�B���7���?��;d�� e~b�����4�cI�6����,���GE��yA�W=`t�=��KL�U�~�Ԛ��l���)Ͼ��F��P�"��	LH�m�O:�B����kf��@�	���P�K�0xL��ӆH����w3�֥���O�_ٖ�y7����dL�>0���ɿ��R���k>d  ̜m�НLj�Ŕn;\(��*E��� ߟ��#^���6��j�u�ê�5�v���M���o	�W���=*�����#������f�6��Fn�UE+ �P^M8}�K��ej'8�U��?�y�\#
��P�]��~�)d�������̨�SH�_�����qYR!չ����;��Z��3���{�H�S]f7�QHd�C�1ʛ��c�O7Ώ ����)�[5�D΀>�87_�O_���̞[��[dm�%JQ�������[�b�a%�٪N���:/�V%�OBU2��nQz
�����K+�:��Hź���}�1�6��e�%pj!�8Ի_֧l�.��D���8�_�car��o�4�o0N�)v�;�x�"���4��i������U��O� a�:)�]��K������͗��r�G�za���{���m6��d�&B���{� �v��@O�W.����mg!Eu�@t�%�*
wT4�#�0����$�$��#�E�t�A���y%�X�#S��M�Ȭ��~x�����R��X��M��F��={V��#�&���4����YUqz����yBpLI,���5�E��67'�ҟ����$e��`�U6���T�1X���V���.|?��9����צR�q'5�`���\g{�B��T��r`���G� ~#fF��-�u*�kqe���2��j�o����gBmÚ���J�-Nw/���L���dϜ,}��L�󂀺ȿ�;U��D�I!��j+P��S��C�\���P���q����������!_NhT���\0`�Uܖϛޤ����1ܠE�Y9���l��+Kk��2l����&�	A���`�,=�ܯ�0��SN5��xҺ�5�?�=-V�C�
��%�K�m�qc���/P��/@~d&���e&�J?�^�	�/��'����7X�W&�r��-�@�an�`ZxQ��҅іan7��]Њ��\��R
65�(��.u�)��UT�ɖ�����`�8�[����C��k���r��,=��w~n��"�>��)SϏ�j�wC�c.i�6�&��Q�� 
�q���;�:�P��0��qᶻ˧�n��
���V̽�)��������N�����]:vr�	�]�k�?���%���cI��g�44��#.�t��.��R����~F������y����R�����O�u4']Ѓ[�LZKe5��{Y�\~���3���#Ե%(2~='������:QDQ�s��"�EtV�L�D��?G˦�T���5��)��QB =�� �LC��o_�N����|��A��z�p�=s7}ҍ?T���i�H��mr�y��;����ٵ�!�&�Ӳ��@��.V�H	�����}�t(<Og�"�S���ߛ7��ܣ,Kf��|�(�L�ʀ���s
;δ�4�!�l���-D��5�)�Z�{E\���}�3�Rm�0��:~LC��@���w6����Y��ʅ�f��`|���|��b���1��A0��Ǘ0b]ٹ?N��ܣΰ��I}���P�B�^�v����ϋ��TiƊ\c�C���Vg ��q&���`��!�&�Q0�˅�0��.��'V��~t����$��E��J0�E0��c�l��O��ر�G��s�3,q�p��+���H�n9C��*!4}���IPͤ��L{�0�}x�W�2�91�t+8@ȃ����%�B3�4�qq-3����bQ�&v`PA�`��
m'�/!��r�r����`,�E�A\��2B��L�*0Н�I��A@�FS�zS9$��<����.����U�x�f;�����x��c�y�1R��V)�h�]��i�3{ڣp���0u�	���������s�_,_:��2-�#��U]����t����@#.��[�-���^��jԥ�%7k@��cD�X�zըIW��PD�����~jN�����E��]kxF'HI�p�J	�Y�dd�f�����b<$�&A���K����z�*�p^�v�fjj�c06/s��� ��HrϘy$h�=x�2	�+T5�w|����m7��v��,8��gi��MeER�s����RM��<����@��pKE^�>G�������#Dl�"�c#�`���p=N�$d��9�ų��a��f_�I~���+i�+8���lY�~J��c�Hcj�˪�:�+Q"p��roV��>��V��&"��L{�E�o�PsU��$=����V�ٵ��RO�wz�_�Z�vCVf
+�B�w6 3Q�"k�*��!�x��`��D��6<��ڭ0�gu�����dV�a*-�=��맀�9���Q��A_�� ys��9`��pσ�D�*7��3�tL�	��E��V-�.6�e=?�\0���C��*�F�@�W_��I�p�{19 w���&ԗ$>��	A����i5�'���w����AXQ��K(��ɜ��������n,D�S�#�"geКvϡ��c��箪/�E��5eO�Z���A�_(Y�7)ԏTh���]���,"�f;(����,�:CF�����v��>=�b�:�cA#�(�zO�}��͡��Jj!��(�6�����ڍ�^��N�u@h�p��zn�gq�B���xb���g_|�8���2�H�V�X|O���٩�Ž� ���t��h��6�	Ƒ!�u =����0���f�������^������%Էz�ϵ���������ɣ�"	�Z�L�
�2J4+�9�kq�dܵ�K��ds?ޠ��&��4*SU��񟱺kn��J�&	\!bRK7�i���:C���]���(
MB�eC�rBX���:��ĵ�������Ы��u�	yq���F~h=�2R��vY���Nqtm����4�7��>��)�|R���Q���LK�G�Ԯ�!D���K���pcSW���lx�^����� (]hm��;s�	��˛�oK|>����IV�'����/���%�;�R�([�\������I��o������9��e�8����=Q�\��<��YuY�݇o������)o�S�'����i��zq%,��j/5W�e�@��?�B���\�<�.M��S���;�}E4��d��Ul��$Iu�� O�k��w��S2Tׅ�	��'?v���.8���V���YhMbC��fs��nz���F��tX1�����.px�κ��ih�J�ȿ��F{�_��^���o�����4��t4NoOP��Ѣ�V,F�k�-sT`i��7�tc ��"�y�Ck!���>�����s���w[�ݑ���a|�k�v /L,�ʂ��Z�C5�\L�;	���H���\2L���jM��э��H���
�#!H>l��&]�m��vMR-�>�dU[\�KfsD�yW�=�z3�3����U��iñ�a={z���pWm0WH/I��H2�_y6�xƪ&E���Q���~L��~�2]Q�E*� �f�Z�P�gG_��@d!�)����08u��M��zP�noRa�HI(�6)�~.��".��U>t3��_\�אT�~�,x'�������(Yc�{t�H����jH�.Cb53�u%Hv��<r���qK"=�nx�Qaܮ�s2v42JL�_ Id��*��MH)9��b��]Χ�g��Zj '�\*�5�p�EC�,��љg�&�C��U	r�[?��#����K���ts�؋?�-��350m!I��[��JX<ʁ��5��q�l��^H����BGE���h��c�f���t�aCt�z��P4�������,�(�4D�b`D+�ړ�։l�%����ja��O&�0�!�L����F�ğ��f�J�8�nԸ�څ�Сި����y]b��(��Ũ�e5�LZ'FY/~J���˻�G�?���p� 3�Ż�q��d��YY����g�ӟ����`�3��S�t0&�d���|;������`{��M�c#�^ୄ|Љ6{QW̆fI��WAˍ����ȯ�/�O�fvGh�������:[g��I�{����X�1ܹ���;�nUg�(F�6�NݘmҞ0@֨�^.�kaB�L�9����2i�ʋ]��]B����.$���\Ld�e�(�ry��B��ю}qk�j>���7��M�yL�-�|�$Z�+�����o�����l�O��a��8����E�6!~M�0����"TPq��`E�8��G��؝�q�.aTԖ�^��ʠ�I��!�e���^.��%����3���ʉR{dn�{�������s���{m>�ǧia� ��3�bm]�Z^g�HJ1�8k1�FT�@؈��gQ�'��K"S��r�Y�HQ�.�k�1�Rz� �mri}p�)s7{��	��"���n�J���`j�W�e�8�����)��%���4ƃM�4TǕq%�#���
"���(iv����]O�P^;��c��WڬG�^��4�0`�)��RF����D��J�>	#�X5�hQ�)�᪸��"-oDēw"s:���*05�x>w����V_$�����y)$�>U���\��UPƏ�<W3�3C�������n8���6�H�o�JAE`]!��y@C|���m`����(�#�����s]#�pH����q�7(�jK���f+u�%)�rJp6Y5�}'Q��Ҏ'؋����ķI�����M��!��/��@f����/]�.O�˛����p%�Nb�Xcv���s$�i LZD�C_�G I����kI�!lR���)Q7*��GN�@s@�"��x�
�>.��+�wXB�|���V���$�_�����c�?z�o����{&n�4�g�C���Ԯ�?�O�7��yUj�7&��s��b��h�R��}!����q?u���iar��7�S_&F�����"�k]s�����䴎	/��*I�M2�|)BB�*j�)�\��R���s���{�]�-�M��`ɬ���ZkvY�2�q�
�����u�jxA��N��E
��� �Y���c��
�3��%�j�7���G�$�·��j�\?�����]͕���m�� �+��Y�9�n~5��Cu
�(���CCM����S�/�˩��㳢�0|k�?Ѫ�W��9i׿,��8�yfT�_���_yy�/ב�L6�s�������j�.�	�rP�2�����5_6�[o�ױYO��@sf�=d��v����<ګgJS"Z��6(�"�Rj����o�e<�*�&!m����uG���h�Dz�������`NDT���C��	���h�I�q�2�a����[}���&,}I����z��0��j.^յAC~��%T#Z?y�{�))�eFP�{�69dP�~�O�|kA�@���§����Յap4�A5�Mr�̴G����W�r�Z��wX��E<rz`��!T�������o"��X/���<<�Q�\u>��86^�Mv����K��I�1��] L��[%�E+tF��[u�t�`�bU�-���T�H��4
F� �!����4L|�@gUJ��rsg�Ԉ�?A��lD%p�ꄋ��4����H��`q �-g��!#k��k����4Ԛ��D�o��U�R��PJ�Z�9�	��[~�)��.��u�{�6�t s��m�>�n��h*��]|pu�Y�(uĵ���x�)���m'�Kө^�ȟ}k����J<ܕg@��I��qw{�{cMW�� ,�9��n�k4*���Eb�ZZ�%3s0��P��:V%p�G��Tc-�d
��M|��(���+��\}5�� Q�Y}�{�&#�~�W�L������J�=鋊C�0�l��2-U�VO�ݡ��9����x��ǄmEw�S���;�]B��0�=�'�7�?G�A宍�9�5Ο�UV��-L
�4#���7 J��i�N�!�Db§<m����༹��ͿG��Ep��2�q�dz(ߓ�7q��S��g�bU�#Qf�\R��b¿i-I9>"W8��y��Ņ�� mO���Q~��J^�.'x :o��O�H�ŕ�Tg����]O� �����gn�q証��pe�n9���¹���ko Ek���z���������"�;�O�@t� ���&j.A��=�J޸�A٥�]�\'���|�a�!����F�E���c����j|�Z�� �/E���Ф��!U�fd����Kf�J"gCI�2S �f$L��~O��N�������)5�wшi$0� ����� t(�N��~v-lS��00>���
��6�0���2��W�I��|��[��`�L3�����ah-�������6�a������wJ�'Q��ht�Ɓ���ȍ�ʹ;x�R�����jY&į�4:zeu��WMY�sP8+��Wͦ@�`�8�/�1G��+A�ر�?���Oʍ(Zkk���!����t-ϣl�����B�ٷ��ӎ�fmIAAz�N��EҤAY\&��y0Lv=^n�0l�j���e�(jf�����X9�h�!Wk=0����h��`a$@��m8��`B�vm*��|��x�2$��7�W5�j���8��_�*�e)K�SO@D�w׊���S_U_�f�����/I�Ԕ�(�c���t�