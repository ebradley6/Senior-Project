��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d้�^��r-�>��s �8������h�Tw#���#/�x%������N+*z�ăZ�4;L�
᨟�P���w��#j�W�iGi���_CPp�I�����9�-����yi*y�k �`��%����\c)��M�wfE�X��G�l�5N�K�6x�S`�^�U*��b	 ���5��G��r>��T�CF>�br�Dtݷ�ǰCD�=����7����Bq�%�(_q�mJYT��U�4R�/��~�/�?��Z~���1"l��X�o��vb��/"������Q</m	����W��
�~�d�K=6܎7��0��h�#��,����[0$M�6�[5sفKjs�/���� E���~z�Rʉ&�>��>�k��g�����_��bM.����i�J�r�� �{�4Q��s�pL�*Vo��Hmv�=�l��	�@��yQ�#S�b<�?� �~	�E�TM������F��+�͗���ve���Z������Y?���Ly��E����B�k�8�It���w���8l�l�F" זm�L_�� ������^���;qⴱ�d^M�k�X���ժt7����������?�Z��p�c9L(���a��M/Z�t
�.��%�A|���B�%-�xDK?;�t�m�D`|i����D����9~�S;0��0�ô˨ "H�tG���z��R��%@�͟��5��#3�U[����Z7�M1�4�W_犙��HA�@�H��p�8�8�����E��Ћ}�+?��C��Y��g8�jJפ&�ofP�긦�~��Z�K	�m�y�,�s�S�ob�6�µ��*��>L��&���YQ��>�aI��ls&sH��K�a~�g^6�Hʁ�����$G�l��R���&��Z}�Y`I��`�m�%�3XD;a�1w�|�:q ��ڳ��
P�z�w����̈́����
3���{ˌ�hl��9�.恖�^�{��Nv �\�zXU�SE�����s�A��U��R�}���vz�il��L�Л����~�>��-T$�=��G�4~��f��/ ����6�uTߋXn�ʜ�T��Gt��U/Ә�L�:!�Vw�
.��EőR���Uym��]�J'��l�¯�tl��u�����(��RGu��6v6 ܗA�k}�2��������{��s�Y&d��#������|	3�UXR������{YY��ȁ�D���t#��8J���M_!>2K2�a�({� x��#��D"��$R��}�����w������U�SZ�Ķ��$�n��^��.Ѥ�X�������AFw��E<�z�2-��pu�=v�1
:�*Xb�A���ۨM��|���Z�RQ��/��+~m`�-Kq#:����W,i�.�ƨ�����Ş"�$׭�8�ž�"�o�e�9`���i9�1��ـ��Zz��4��ƣ_��U��]���a�����m���a��CWuB�w��D'�`�/�~G^�8v�u��Fdxx���0���~J2Ioq�@Nc�]�6�1LpB��fy̝��IfK���M�}�*������K@<�7C'��?-���yY�Z"Y���8��<�d�c�y��>%ȭ�zF��.4Y㼔"��Z��} �Z=L�mJǭ5r������ �¡���,��~��O��Ž���6�t�x �2�h/�M�/���R����J:<�-�Ye_~QEF��A���$բcf�� z����<D��y�A��Bg�7f�c���nB��=����V��(tM&�����Qϴ��a��DR����ԓ��5�459nl#g٫H��	6Qr\>�ɟ
����o����x�����~E��vOy���� �l���
�P�onIr��G,��ͺsܼ��/�h#��#P$8�C���j�r�%Vl�-U�1<����,%����傲��@�迧���_8�V5�v0Ѩ��:+T�c��R$�g���*k��ŷu�u��K]�*��}3>���R^a RD����	\�Y5-��e�=ڬJS�`E���k/e_�֕31\o2� ��ǚ�Da�!��ärh�*tդ��	K�ó�ͩ�cOCE�Bxu�d��y'R���T���2��a)��^�����Ck�(�@���6�gq���69Mv��=��QL�UD(��Y��,��k
���+���R�iၧ|����ħ�(3�K"�^PE�K��y_Y����X\�A:�	ϔ�\�O����B�X�u���CQ�V�f,�0ZEz��Ԟ,� }��s�b"k�ʄCu��.�ye��i�O����n���4Ҫ}w��Q�m��1����R�WJD��G�cQĦ{J! {]�xkjgE]W�&n��,�Ye���y�n�=�kś��?���=c��DS�.%���H�ݺ�_6R�'�#/zzl���D����a�Mwv<D�5�����A1_ʘ����-�� �ܿUY�E{���v�̥MAFcL�L�8p���͕�iU�hIB�fH�� f��I� �bM�+W�͏��LTe��qM��r��)�[xΛ�@��H��\p憎�)8.�Ŗ��`5E�O���D>�П���� '@�a����n_S��U�}�U��v��k�5��[�;�Ͱ�FLN��n�9�\xݫ;S�/6t�[ �7����-�6��;!�m%E��ЙU�Q�P���u�~�W'O�F+<��';�3H�>�IF������*��R���k��c�pC�t���֦����_��i�V��Ü>�i���!�Y|���/��@3�E:�ə5�耰�O�v�:��������b�j� %^�2�v�,=�f������V�="ׇ0��U=*���*�x���q�2O�B�'$�!$�E1�h ����J�J�Gq,!J@G|v��-K��3�F
n�{�dP7�BH�\W݃�J<�K���/+,h#I�#(�l�LO���Qz�� ����>-^wT��W�uc'����m��
�Hq}�^�1�������e���06�����o�P$)�i�Z�"�1��������š�Z�֏`eѓp������?��hW)�u+��e6�q����w����;�U�K"力~%�����b�݈��C�%�&���/�-͐5^ ٟ��7�f^���0g�5��څ3��dBh��iSF �B��)A�|/E(h�Z��=�ɮ�e�^t曞��e�:Ȏ�k��h�Ȑ�b��?���B�:w�W����ΰ�r�u�S��).�����T�����M��p	���S���U��Xv ֝����h��.��vn��4{�y�o�㢍BD����':����g4옻��{wSQl�e�IMS��Ap��U#�2���ⷦzB�6s q���8tS�b��Ѡ.$ʡj(�-��|6Wu-�����u�!�Y?Ӓ����"�9G֤@����W��Z��3g�4����:�o���j��a�T�����w�G� ��e�C��G�n2��0��M��!�i���O����[��
L� ��<���i8�`��������*�XXZ�NS!�8'E���k-�jy.hIݗ��o!L3����_
��7Ì��}�W����Kd<����D�k�e x�ì/�,'�zq�|����ĨVӏ���^�i�`�v�_�&+X�S�{��T.��A��[�f�$�=(<mS��=��p�o�-9���cT1
�	:y���E��D���Rm\�_��L�x6��g��5�4��F�0�t���t�q�\<t���גQp�h�E�.��}U�gY~����k|29�a�S%ꨨ�=�2� 2�z)Pʦ}��9k��"dj������N��&��kظ!oz��՛��g@��j�!�5�W|�R�䒁8������Bأ1�ͻ%�������^��W���᯲�O��l�doM��Yva9��E�Ф�H�Cر�bW�_��gX���2�3�N���>K˹k�p���3*�xr*��8�����L�e�ڐ��s���@`/������1#>_�x
���D����C<��{��{=� ����̋KnJ�ېr�'�$�?b)+T_���6��a�[B�}E����D�3�E6�r�����j���̓��q ����o��"�Ǌ����{$X j��SSR)�|��~n�7z�f-G�1:�X=�N��-�o!����c(3����]�Al��4cD�r��`��]J���;x��/�=!��[[Mq:��.�S]�ᾚ)_�5tݒ���{QX���J���Ē��ܒ��܄����h��c<8Ɩ��HC��z�9w�����	Ҵ��F�κ�G�~���=��B��3�~�^�X*�g������\��k��TnǦ�he��nm#�B�юh�u���T/��S,na�� ���U�W����/O1r^���{�|
�G�U�R��������c�/3LT  ���MO�2���YqѴ<Q�iT%&ҝ����`��w��=E֯�S)�<gN���"�L��'ɟ�`}2�N�u5�t�P� T:)�5��mM�\o�����Sđk��~D�d.�� c� U2��r�#6�LYČ��sel�:c���`	ep����	G��ګ���b�Ut{ďN�Y5����ҭn�Y)��x������l��U������vT'7;{����s�	����kB�ȓ/BX�w��F�0��<�SrUBUF� ��<8ǟ�N;�O��qnbZ��K�4 �zX��r�F�f���T5|����U�Ę��+�V��DOL o�c�]ٽ���7h���fzB��	Q�����f�r	
�N?C//���`���C����� e?�@�`��"�]�����]�UA�ES��O�^���1NLX+3���4��gJZ��M�{|hj�N�h]�uVE���U"&XN#�wƄr�5�ӥV�R¤vS�5��[��ɍqO�d.��L��>�n�z,�DWY/fx[�a�$���E&%��
��
�	������J-��v���B�*$5�z3�
�ԿD����ţ�5�Y��U+��bR�4C|�b�C{8�H���_��JG�%�����mA�`�e�Mmiɼ<��_���B�\q s���~tO����0߿� �+P�z�ǌySXI4G,�% ƒK�m��������r�D�\߈�sv�0�
������T��Hl���s�
f��䘱���?"Y����C��6E����L���� ��I���ˬ]Q�6�	g�d�j�y�ʰ�	^?7!s4����ρ"�@|X�u����K��p�(�U�2Y/*��}ي%F�����q�Y�+��Dp���Y8�GE�2稓B���B��,9R%�Zn��<e�&v�}}���S�V&�J�SfXR,��<O=�r*�Z��f�sS�=��˾:��`�΃��(�L����w�	������w�<�;��K	�~���t����p3�Ŏp�{F�g={��Le�"���Fհ()��Z��G˛�u�]*H!�d���=I��+ac1��_8��|ӑ���;�T�Q�;1�6uq4l�U��J�E��������ty
����{t��m"s�u���Hؕ�4�q�XR�n��h��X��h.�����J�5G��J��R��?��j�o+�����g�Ċ�<���R���i�>�!I@W6O�kMP�I�WQ)��f;�����rm;�V��>@;׏�":֫� ��G���U�H<�bYN������jP����6�J`V��ɤr��~����)���O�U5%w�?ֺ�Q}���Ż'8�E>��^�!��{L5N{���-?�R$��_�|���B�L\�@��y�H��Ö��Vm8(�����%y������}�	o*��J��9c�����a�r��zS���s���l#�����Y�c���s�J
�(�(�<������Aꘂ)�.���%�݌<�V��Ag��9v
�'2��@>�EP���E.�TQ���CM"�4F�Y��b�[���y��ju��������e�4{���e�μ�uO��tB�uss�T0.k�Hh6�xW��s�Q5Blf�����ft�I�����K�� -x4�5Xv���R��O��.��瀶𛖞[���g3���EP<n�)o��B>C]�O5��F_�q�Y�r8�n_�7�N|%�ĥ8�����c�Vh�@�c��� �u!����/ز3ߋBʣX$�3$�JK�_��s��zI�O~)�V<(��>�b���D�z��&�W*���ŭD�1���#�
`�ڴ\��sW#e�?�T��7���k�s���,6
�'�'�9�[ąGaVޡ��_T2}�Ư�z1�C����_J��m9�ψ���v'	�xiW+�Գ*be�"��v;�k[�H�r
��Ǚ�A�-j��\���H���뭑�΍�1KY�?��Si+N(���G#OS@�8���"��D���d�_�|
BD�ٽK�D���cyw��
>���1z��
i�x��K�뽐*}�������M2�l<|n�72�3^�`�W�#P�y��f՞ �� ��v�U!Ő�u�U�Fh��+��A�Hiƒ�!���N\ų��u~v.2FɯrQqV��'�m¡%�4O��@f`A'i������r�l��|N���9|�/̆���\7�fY�?Tn����_�����a�d��o�q����{{��W����
�pL�3)��N�o]���������������1����%xnN�e��g-���t��&`�nAV��-ݎ2��G#�64�W��z�0��q,p�5�M>^r�z�d*��=e�S��'=�Y-41-�>�h�#�I/�`���=<ڥ	��F?�w-�b
&�}u06�RS�(}E���U���?�?}��z3L�e��ˬ��wEU�"y��G�>�>�Ώ�דI˼�Vqʍ����'.Z��U&����d���ͿR��ǰ��	M���%����@I<�梤�]���MZ$5��Ff�6pgGlMJ�}{��\�h�EL~�����n�x���IA��$@?H��H���E�W^�uҪ�&ւx���Xq�ߨ�����EI�`Z�1���JB�`:�ZI`�G�84��#�Ftf��7���&����Q�f�4�L���!G�7b55:����G���k�r�k!�j�Hf���)�W�~h�SHξ��D���(SZg9�"9]x)���w�d�ߴ��|J�?˙���BQ�[��Z���~�X�!��5�#�a�i�����c�	�&j	�!�r�#b3Vtޓ�9�0ǌS�p]%nT��X\LU7@�i���A�K$����4��!i_�*��f7 ""r�����C3�	<�e����Sz��ҍc�	2�م���P�8^�B����['_J��ْx�W,��'e���I��cmvh�Y!:���c����5\��Ĉ�1w��*-�}���Բ�I�A��l��pj4
t�QmP��c��XZ�$٤\`�yÅ��Mk�N�4�nL>M�����<�]�/��6.���jT�6�,}�SY���F�a
q�����
��C϶��f)ekN�Y������CL�?7��eMm����6��;��k;�Ad%/L�	�K���-�.�ה���Gj�MC8yP�V����X����#���`2���ڞi}�-�f�O�Ҽ{�t��@��h-$��YZ��ɴ��s$�Z|��Oi)Ά	�$�|�o��n�����ɸ;���p]��d��GsM�蕮�&���쑨��O?퀗EI�BvA܅�TzVL�-ťح A��gv� +4���`H�k�^Q��ĈM�$��_?��qwT����Ė�A	�pn�;΂8y�!1�Aq�4��g������W�֟���MP`�Cc��%��N�`-C��L�3�o�e�J�}�+����!IY��[�A�j�z��/ݡL6������t�xspX��	�W��YI �����?���(Q����f��mD�]n�y��6t9����Y1��yd�����w�ZV�Rd{�u��J��x,�e��>�S�z�X%t�$49m"˙���O�z�i��q[�R8>�سk��myd����q�pg�C�f�8ֶ	t�B��BS�� EBI�W��c���N����2Q.��%D����h"��S<��"���vZ|���I�*�%. ��ۙ쓕ۺ%���gS �̣'��_�ey)e��� S�2p���~�na"y�A�Z��^�,>|"��a���d
�'{��Wm�� �z�����г",m�-�����*my?J���E<�Td*&��J|�i,�wP�À~�;ң�ѩ�[�l��k���0�N}}�!�sbK5ߍ�Wawx�\��z>�8��Hl�K�o��1�9��/�u�K��K���X�עn��c�3.����/G�7!A�|:��Z,�� �ĝ-��Mmp�+2P�l��N��60�uy���$4����i�퀑}Os��]G�X�6�(�#�7!�m��1��[����爵���I�$��������V�E�)�sJ�(��w�w����C�a��$�1ۥ�7QwʣN��͈T�d;	fJ/*UY�x�]�����D?���5���[�sfL��v�-�}����d�%zD��O��oS$�Ё�(���{�C�;����i>�nͧjY汝,�0�lK�tN��4�:�TȨf��B�;�f0��$�X�t�]�����?i��,
��F������.
Ҭ��7 �F>zL����vP"ŬZ�5�sI����y���!�{- Wg(��i��ðH����X��:�m�:y�0���3s�H��$� ����yF�nm�ۣ���!cJ.�҃G�V0����ઇ<�����E�W��`�X�5�������g�TʂG)P��6P�qw�h����Wʒa��n L��CaQy�Xj�����:g�l��]?�s���j/@o������3������^�iD��ݮ�o�|��\,tQ���E��۫�G4�8=֑>6�ba�a��o��X�����=g9J�>'�1�4SM��i�����	��{�ۜ+^d��4}������n2�F�uW"������2�ge�@��0%Ĝ�xU�_1\�B/�G���6;��������u�4&<E�Z����:23��փS,Cd�K�����ٓ{� ��L�`*��%���0O]|�X��,��D]�l7_�qoXӣ`G5h��β8�\��V��n���qW,��[&,��Ӱ�t���"��E}Pup'+rK���75�3�ʌ�G�o�Mk�g�,^Q�@"���Ze[�RiM P���>h�V��qgB��Z�R_5G�M�,��
1��Kʁߞ���f+�v��&i��YM�� �AT��gET�����Ӹ�	�t����ݍCq���sS� �]�E}2|1:3͇*�&+����NF�W�	W�fN�;����p`e�&��O�3,ٸ�	��b�ff� �>����i'�X�n��o�"Fs@v�]�WY���p����I���܏Coc]?�X�����4���R���:}M��3j������4���� ��ݐ�PY��(8�Rӕ<4�f��?J ���o=4�#������}3����2�_ܿ�w��n���|=է�]c,��-��r�R(UO�_B���I�J�:44ή@聠����v<��H���YIE�1���?޸&Uޙ�ZJ�9��]>Z�����4����-Y��{���Py�j�A�[IU)������[:
�Dc���d9����H�ҟK'L��\�����k��0Ҵ��9�y~��Q}*��]p�lrt�f`l�ޓv�4z�E:���(�_�g��&�F�H���gF�>�PA��Ѫ�� ��~�4��&mW�A��2����˓��$ܹl��Q�ߩ��h��ڢ-�{[���V.Q��L�}����6�U3XNX�����;�� ��c~���!m��}�l��C�tQ�LfP9�O��G�$�Ƥ���>=�
4m���n/�nŜ������P�RJ�5-�p8<�b�Jg�WQP_?�y�MI���u����UGT��^t"]�8�P_j�w�<�W�Z��Oz���r1q�e�,/���^�Y��@�ί�W~]����<����@�t�E~����ɬ���!� |:ϥ�@nHмGo�IiX�ו�`X0m�?8<o�,��N-|���l(}�H�Ǖ+��A��©+������$>kц	���O<�qg����C�f�Z�E;��ɡ�A����3��-�P�T5��Ш�pv�K�V{Y|ڸ�.�_����)��
��8KO8��
k݁�ĬH��A�_D�í`�?g�l�U<gڷ��c��r� �q�))~�z'r�#�5��~4��Ռ6�O�|>� ������v-{HD���Wq�Ν��Vتf��w
'ύN������5+<. ��&P�S�����:�mR����1�D�[[#��Ov���Y��nm��Q�ʭ yF%��y�Oc~������:5`K;u��ҫ+�ko�gƬ`I%���dhs�&T�.��h�4Ax�FY�����]����Ȱ@
�i��9	Ռ":�.�bg������r�B�xqYbGj�� FN���fUkV��_=E��?�j�a�z�k�-�7D�+�TԖ����Qt=D;p���L;V�Y�'��A�lv;��z�s��LZ3��������� *�ij*�'�]��6��V�i�t�iE�Ύ<T�G9�~�`�5�o]�A�1�9{J������8!�Xh>N�;˱�l�@	2䛮���YD�ɧ&��=�C䅹���z�g��I.r�-�LZߕ"Pf^VV�_}��������;(����k�G���o�����;���e�>Kќ_����A]���ǌZd~�b���7��~�uP��x�آujŌf�� ��F���fDg���(,t��!$l2`�(XL��XU��]�q�|�q#��ze��6o�W|n�u�pi�r�A>]�g'33h����q������{��׳$k��"̞L�	�����7��� �@��!���O��M�ܑa"��������+:h�[�͛IΖt�؀��۸[X58t6I�0~n's9�w���aS+�������%r����jr�NEb���g;ؽ&S���#������̂1�5��n�&��B���c?O�>�?!��N(�� +�����dC��؂v�.��'����aU���/Q�����_��A�����2���}ycz��@��c�Y��WϚ��(�\�HR�������h=W[�J��!�}��������oc௩^�z�*����k���Q^�wfP�6A���g��O�êJzFy	=G6���(7�L֙<�V�k(���	���<烸��e��h�X#r�,J�u��w� q>��De�_	q?��)/�hV��"�N�4�4>uc�-k@Lۭ�k��3/wmLT��%ޜg<I�H��\�t6����y�8��Ȯw䤬8����6��R��0�o��VDm��ߕܚ���"�+�˨t�qb�u1�T&�*GG̀Fw=����a��.�]h���F����\���ހ�틓QD���]U}�@�ה�6rS�UӺ.XQ�!��WJ�QkzA�
nO��qR�m�I���ߢ���>N�.����k����Pȇl�je����k5k����ߌ]]�c�x���ݪ#��Ѯ=��q/]"��w��F7@B-b�W� %d��|a��$E4@�n3D4�i9Z�|]�c4�E���a�ۍ@R���B5G�"�=��'x+� 7�_a���M��А�
9�O�.p�h���=Tژ� �6F��c��2bY�`��!���6��}՚�p7}��j�I:�����n�,q�x�$��\D���E�����!�����¢�a������u��Dz״�KW�g2rªʕ�3��U: ��	�ųfl]��:x?��^ăA�~��f�F�7��]�A(a�ùV?�ś5�u���J���>eJ(�U�v�[�Y|%��S��z��P`���PH4���B��>��ݴ(V�+�^fPբ�wt�aeW�2��P��⯞���k��� !��^�
���X]�1U�^�QA��4��I�p�Od�Hй�bȖAT7�P%�#7��z�}�^��Vg�}��)c������d���J�,�~��ea-I�y�u��^$ݚE"/W�wo���DK}�7�L3���g���ExuC�'}�gG��:�(b �l�L�Xz�뿙�=�;%(ʖ���,(ۅ��)��J�W��nxO��aU��~���v�'��w+U�t�	`C����,�إUm��b#���@^q�NĐ�����+9}����%������>�E;6��h&i��D+V�wn�%k"5��~2�1BTc�&20��|��O�	�<D�?���=�%[�ֽ�R�+�Z�2\�� ��x���Ӄ�Bh���*��O��ΛW�:>�p���Z��wT�5kc#�7���8#�k2��
�C�W�����g?���?�L��*h��|�p�Ǭ.~������Ĉ�g�q�]�J_� iW�FXA��br0W{%������2���<�5Ru���}��T�<A}��R�����ξ��8U0��sOw{J/8Z�����|�x0�C���/�������A���6]�m>ST�غo.>��}�$�ֆ>p g�jiW-���>�yp�������=�x�]����YE�x�m2LM�q�HΧ������S�A��W����K;} ������-�y��[��{��d�*��t�L?�<��+4:�b{u)���klU�m�%��˭�G��=�nx�q�^�*��Y�Ѣ �~>��#g4���I'�U&�ҽ%�-�ȟ��X�g!<�@W6���nRg����}��u��!�8w4ڹ\��3��([0��b���(qp��j@m�1�졓Gi��U�mÃ���֧��H9�Wj�Y(��i���p .��c*�@\��f���b��DB�U��VP��S\�|�@f�'U�g�����ż�+�r�1o\�4�Ɔ��Q9���U�H��Ӝ�B�)��4���]�|�����Q5�Oߔ
!�^�����[>B�S�p��U���0w��j#�
���+!�9 W�?8pk��9�C1ݠ�0���\v��ě�Z-hڗ��ƼX��gz+�w�@`������d��2X�`΁����\��31��/����Rj�����K!���	�v1.��Ubי7��@磻5�A���&߉�:��]�Ԯ��	τ�۱9����|�b)�W;ᾳ �H�E�rm]]/e��63!lWc Ɲ��2EI���"�KZl�^��3'�v:�LHZIA/�  ��Z�,`v�C�$�C�,D����*c)\[?��oGC;��
�~K�G�ڝ]��G�CX������G��m�Em2�\�X��-�ݓ����+jEo�I�AkZU�];+m�� ��F~~�4�U�Sb��N�xM˥Թ{��q�@��U�\l�&>"�)��u�QX0(��]O����
H���N�8��!�?���H��i	{bj��U~��C�%H\mD��f�g�\�o`(�qm(oU��*�@��Q�ӽ/*N����ʼ��[6H/<����n���/h\�KA_�6%�c)B��!��"���z��G�Pށ�����%����:��L�w���T��уԼ%���'}�QҸ;+�ә)1P���n��cO����N^�tΰ�<����7~u"�.��&;["76�$��Գ�wp0��p��?mO QƧ@�##��hO��7*�u,���%=#��f�kM�q N�j�]B]�lm	�cW�v�?4O(�ּ0~����5��C��h7���'��U�f_��)�8yj4���6�P����c�ߠ�Re���� �,��l>]��������I��eeUm_1�Dޥ�{�Q������'�t.	���"av���A�lR�:�?����]P��mmV��������?^FՌX�c�5�Ӈy;�V�;�/�w��f�����~=�.Ԅ]'s8�6�o���}$��A�T@*s�7e��5��+e*4�O�]�`Vy�����E�&�#���$q��A���>��d]g�&���1ᐥ�(���- ��x��"���V.^ǪUW�)ܿ����=a�������9r�(���7�����"I\V	UV\��MH�=�'fm�$�������ܵd�N�E�\VoWVY�!u���5���i��t�{4̓Y��� ��i2��^?����ج�0)1�+`�(|a��wZ�+���#������1���m�`D�j6�����O��X,2A�۰~��Uw������.[��a[g�(����d���֨����J�Ï ��@Y�wAp��};6X�3=4U�F@}K��(�{o�t�f6֓��s�;,B��k��km��Z���V�*�5��$!��H�G����<�%���AB��pC���p�0p��%\��g�,�B}���ͤn2�@��H;�6@Up>�(Ĩ)��f��ӣ0 �&뒡7$Ku�W����+�2���4�_��5�\�s��^�
t� ��A�0ߨUг�X5{��\��3�bo�m�-����P�"A]���L�qs�/���fb�_2R������X�M6�wZvF�8B��ni�!�-B���T���xf<���*���2�w���Y�
C�x�u��d뾷_�3�?v"���o����^e�}/ԑ�$3&1��*y0O�'�f��$9<���O��F����v��� W�V�u�l�^�n[-(pg��W�X��ODe�k��X�j�q��J����U��ج#]�!-d��W��M�0���u�r諬�D����5�m�@�Y�K� dF�0��	J��>��e��pt2���0�4"�_��b������k"?%,��K�+�R,�Vd_�N�ݼF�������R�"?B(���O߅h%+�DtX5vD�t��wBr?�V���w�$�h��ǉ{K6*��9�b±�+$��ł�.o���)��B��r�.}����;���Ӭb3��#��&��H�x{��ܷ�w�����`c�%�\�v�_b�j�w����i��J���[}�]W �����7*�Dx����>�r�'r�L ��JV��&hA_�W*��J��Y�Xq�e��r��^ǹP��Ӗ�=��m��X]z��M�6�8,����] 6��DZN���F���7̋
$�{��K"�/�
=E6�:��C��uۮ:����G�*���9՞����VF����M�ij��7ީ�M�W�e�_'
�Ś9d���I��e`j��4������[$���N���fF���M�����LZb�$��O'���2�P�.��+0=���&a:zG1uDؙ��"�a�\���QV6���$��|>����	�%3�X�����X�R/!%��8P
�(����1�Ў���c�BB�2`S�:KM�We8#xV�/��;�Qٜՙ��ٸr@E��A���}m-��|�͐[lc��Y�{�ᎷW��Tf�qC;ǝ#��a��[�?F�y��$d�s�I)!;^�N�S4���I�7AI� :���g���d���3�����'�=I���R�ð\�L�(A��/��lj���h3pFϙ-'�P����t�P�b��X�Q�$�BT���#��M�RlR5(���w7���ћ����%�7�y�WF��+α~�m��Kt���K�.�JE�!��f�!��Id"��KfԶ��?�E�wR��G,�[v Kq�jL�
�i�.�\�������d�ב�� �f�r��]��"r��_�	P�Ը]�|����*:�K���)�4R5&�"RS  �+�p�R�v���}I�!��!k�g#��ڇ:/$֠h`m� Z�����e��m�q�W�����V4p�}ge����H�Ȼ5V�ːC����?���Y譳��3xn�E��&i<�&಼����A�Gx7A�:3~�H9l�پ���P-��	��4�R�]��o�\iBlx�ݗ/X�y��R~�5��拳���=U��$S�@��a`�hx׬�o�~���7'��G8�H}��B��Fxڕ���z,(*_���t>8 ���{�V���<&Dx��$�g���ot���cَR=E?����9�tCz8!��u�7ajfo�O�p��NA U�nd(����.X��|R�5��?��6r�� } r�q��QN�wz�y~h��SG���l�xE�b@y��w����Yr�@g�%�d~�pu�f�� ���#$h�U�r���	�+7�X�ӵ�D�P��9�l��ެ�lV^{�h8���t{3P��������e�<7����`�K�2��- -����<��#�{�?����O�!�X�p�F2U��Bw"<<��;����<���B��AM��L#ԍ�v�娊qP��s�������vEM׌}���Ҕz�Jf��1�,~:�#�n7{k!l���\	[����E
�<:���b��L��'5�XiU�f�T��Kz���L|t��s�7�����3���m�cw��wn�b��-A�ɢ�>�up�͋��lZ��*{v�9շd�'S6J��Ã�؃���������2P��}GS�1�=���Ƴ�#z�Z���;��	k��!��P�*�7�c⸇MƃR���5'�+_��/�9�4vD���A+�({t��A���'6�T��ے���4���@��;i;\=YYsI����M��
��P�������B��F)DF!1�"�&F�w�G�l��+(R�Uߔ`�|��)o�m�V��>���Ex�_@�0�)Z�b#��[u��B�rwB�.O�慭�K�.#��]�w��:�	)�O�W>̀$s��w�� �������r��8��v��_����N��XL�����c �ٓ$X�,|����迤y�k U�����e��P�lTc.��Hޱ]�_Hg�����q�f���Kh�.f�,��r5O���+ ����?V���,��s#�L�hq~F��Ja+� 7~ʂSt�MF�Н��D������|	�	�oZ�~�p��W*/Y���;c7���sM�!��oA~=u�j�!	2�5[*�T��v�])�/\G��R���>T�U?�p�'//����j�2l���
�ӹr6����F����u<`^V�B�r[i�3n�\�T�?�n�������%RXY}f�0�:��� �e�@�1s��S�-d�S_{7��8����GF�����L4 }3��B��G��(�z��
[j��Ju�h�i�x�vq�����,(v�	X�����u���8���2ǁ�P�3�����z��Q�̾�a�0'�d%O-��Z�Bf��!��C[o�z�!���ĹgҶPz7d;�0<4??���Z��Y���J��ma�E�p�����t��ʫ{�U��d��Ke���Y�m�������H�N���2y�e��Y�4��Q�})+�Ҫ�峇S�уm����2��A)�k��
7�(���8���v�-�s;�C������}JG�K]A/��LDq�� E��B�m��`����j˹jDlf�z�9��S6�'�R5M ��<R���6������\ ];uM&�V��dxV:��l.E+bA(�y���[-iߟ��$���FO5��Ap�:.M����[U��f�0}x�� r�*�ș�:P?���	��]aS�1d @�	��o�Fb�4����4j#QdW��*,.���醆���w���u�a�y'>�qJY���!C��Zt�j��77P@j]1zC~Ϥ�ߝVR��Q�m��;�$:�.zD�|�XTA��2���mn�W��5���ҹ�S�`	ϗr�-���W�E��;��(p���itU��}9�GŦ�m�	2X�����c+�BX}�<P��2�g��-~�E�Z٪�A���?�7p��?�m?2��f��^��nJ�b	�xj���>Dl^O����v�%��G���w�]�J�gx�k�n�*Y>#t�^t�p�r��U�6@!%�Q?G�Lvx����T���FZ���Γ�˽�s�y 4�v�%Ih�٢�Yë��m�1k	�E����M��{瘏zq�',M��'̀�w|&��o�j��e�E���fS��rJ�$ݬ�.1�G!@l?�%��B��>k]�ubW��#�����pi� b�����kF��(�-�9 D���!�K�4-U��]=��� �ߒ�����89�
v����M�SD�sމ-�(k*�2��
�n�S2����7��经&�E���v�
�Ub{���
>��h��YR�F�?������!�5���v6�X�֖Z�@�B��ƂCjд=�������~�<颃	��!�.�Wf�rŜ��}z4�ۡ���m%'������v�.kW��{̀��>�H���x����5ŷۼXp|akNW;ē�`p%�Y����$[��1dYQn	�F9,H��_�Ư>vB�52��r�G�g��J���l2�������Z��#U��X��n�T�n%�<���XX��?�3b9ey�Fx�I��jB�|c@<��7����{2\��d��2���*O5pQI(��Ѩ;����LwA�%�����b$ޛ��ZG��p����:�0��9���+學����qܥ��щ�uB�P�̨㊹�d�w�=�7� գ��=��+'ek�V ���cO�T��x?e����JV�d��,"M��Z����#)Ǐ?����x�f0����*�9�'���v�Bu�r	C.˯��n��mӎS�����0n�
�~f��W���[�թyx�	�A]��ر���);�9~�N�I�p���n_�g��$���G�����UL��c�e1�a��5���kq��2�d4���<��<�h���Z��v��x�LO��@�3y�	4�N�(�so����/�L6ġ���,�ʕ�gA�����NT���]���"�㠜1���ϊ����T�Я�����l�2� ���W���r�t�; ���Qsy�U�U�xǿ��<UU�5���r�6E�o<I��G[/5
b�譊����-�1���H N�v�4)��	���x���j��ջ]^��)d��W�ĥ�p�r�����wv~��X�m�8�jΰ[�{ѝC���oXkR�����W�r��w�;F3I;|m͈����<�AX��ߍ���d�c����Цe?�u4�I��4��Ǡ��S '���m@@:�q��m8;�m��\T�;�=���<:���aOcY(�=�Y���NT)��nD��vӊf���/,�_�&�qO&
Ԩ.����-߃�3�x��C�D.)wA�9.��	o)�BQ���6_�������ĕe�	Hc�^�g�&��u��(~@�=��හ��N&��I�2���BE.�4:�V�tTf7+��]��A�O�k�;\�K��q͐��/h0���G�y�yt�P�������׾��6��'���pC�g�9���!�Q8����&L��RG�*p-h�Ƥ�|Lf��N��IԆ�����j0��_���E�%b�{�Lo�Nē�O��ߋ���c�tOa���)e�`
�.�޽��Y�]#D)�?9�H^�RDF��
)��h�IԠ\ek�	&6'	pc��J�(r���\}*ؿ�����L��Ai s�]([=Ec+�؁���WŇ��t���$�5�KQ](�J��e;ά͕�}��<o�2�8���F� �1��<��o(_U���Ь(ljxPP��Eפ�F���aϞk1e�i���D�y��$XԌ}��ڄ�`P�9���;R^ǤDtn�q9�t�]��\�tx�z�q���vr�6gpB��!��~8�Z&�7��'1ge�<C �7jB��u�St)v�D@M���]��.ݳ�
�!9u�q��F�n���p�P����~6�1&н���()y��,�����+Hm�9.7U���)Gd
Go�5$�3p����m�OT�O�� �Gvdb^;�"���JZ`M� �GvK��U\�FT�q����:�C��HY��րإV�f���ഒ�G��t�o��p���R�,Q����K��ɫ�-�{����=���Z�;��X:=��hE^Me�uf�b3��*o��Im c��kNo�Kpit_�Wp���9������5�M�/^/YW��̗^X��l-��������D�PXl���J���v�	7�cZ;��Zu3G�F� � C���R�K���b|�%\x��o�>Y�RZ�ʄZ��q�o%|��%���K���	T_ZI�b��w����.�w��F�{??���D�������v0�]�X@����Bs�����c��������mg�>׊+�ʣ����̊���ٮ������{ِ����	m7������2��镻��3s����U����2in�2FZ8AL��͆�ǀz �h�Y�t���`�f����,���&T_*�ְ�C$'ٞm�����j�C ~�'�lD�[�7!,�{+&U(�OI������5�1}�C+R��l�r�;���}s�BO/Y���_�*�ʢ���+�w?����~7u!�Wf[& M�n*�&�6��}��nQĜ�k6���k^�
Ogmqh;��9ؒ��$�����٪S��z'��m���~<|��:���hGP��fܺ����F��%��B2;i�_6Yk�嘔_���� ��2�[����k1���/�*��B�8��;Ƚ�w]�^��X���AȘWs�NS�r��;��R����5�q7�2I[o_X'J��p��?r'��DD�30��"������\f��U3M�Z2�r�2�gQ����^�*����Qz��P�s�ć�6�����}�[ ,���
(m��UV�S��7|�xM��F���&B���iVQ/�6C�JiM���w����q3x��8P*�k��1��X�ň><�i_t�����
���oĮ8��AX{�~X�c����/D�w�zL���>�kI��M�#�$y�y���<��%�͍���Z�v]��{���c�_�0����Ģ�g��N�~�k>wcG�/����z-C�5�Ğ�r~ԸkN'x�w��
jfQ�9�4�,1D`ʍ���&��u��hj� �V�.��DA�w�h����C���*��i�֓N_7ĺ��6-�PHh��?��w��^�f������'��(��'��x�;�.��+"%���r������/x���V,��`���H��lta:���ǔ�$�������r��B;�sw��q�j���~xQ��2xe��a|g�<�9�2���.�V�߸��(a�(���-N�V��L�f#T���!��<�k�n��3s�٢�d�7���1�K"}C��Թ�>�鈽:KT��!���,����0��,�S��/�iϰ��m�M8������#�p�乒Ṣ��@�R7*��}��jh�}^�/A@f�M<u\LE���)����K� v�����޿������a�;/�O�\bӫe�o.i	�JiL�10�Wh���e�	�-^)����YM��
����� ���+�e^�����CuES^pII�ˍfN�Fr�˪=4yy+N���i5\sQ9v_D8*����.W�F����o��sR�� =�nT��y��,�
14��O<� �r��k��{��#��t�WoiđW�P#�(C�pM�ݙb)@mnl�=j���@M���۪�{��z���-}(l�	�_oB;[�T/q����IsՖ^u�%�5�%]&�3���o�>�8�����&� �!t-�p�k��2�n��\�ܧo��A���ùM��	�Yz��:��8=
���vV�A�����0w�%��k��_�6=��Ws��@�1TP�u92�ڻ��y���>N�����r��*������{M��S2�6����ֻ�Q�����	����u����8ЁH���Zk�޶{�sNZ\A�>� Su�D���L�	W�TT��L�_q�#���@I޺,�������pU)sn(���\/7�������mR��*�=x�I��ۣsQ�o�T'tҩ�3O�q�b`[���w��\ �3nm�uq�R��c�Y���h�z�i�}��������&M��->NG���)�@���XQ�*V!]�|[Mj
�L%?䨪�bʇV[<Ḽ̊0J�5X�*�>�\��jv3�Us|�������X��Tk�S#��?i�^��>��� A�Vޅ�IׯO�Č*%�ф�>�����$S�!�=�a�`@~��yZ�u"F�5�9�6��!�rD�/y�s�zg���M�eQ��%Mˎ������'*F��r���cy3��o ]�|	i<���\^��	��jV�"�]O;q�$�N��vB�xF_A���2,/[S<?�s �:�����x��&�J��Ca��}R�v�[��K�0�g���q{4׶�\m�w��~� i#�e\N�A�jP� O;���&�*�N�֕�/�������%8{`h��&5��H���n���r>4�\�C�����Af��4fC�ĝ���k���&�A��oS>�ʻ�����su����WWkӟP%{��a4��9�x%�l���c<�������-��,c����7��-~ ���Q{�\�*�>U�>�m7��� +Cꣽ�T�A�j��fV��2�+���.�c��:��� ���q��_��c�o=ks�f8����g���e��!ЖA S���fy)��ս���ە]��hB�f{w������+8��G�P��,F�ov1��Af��Ⱦ�/_��4���.�������}�U�E��e�b�ȥ�h��L��'m[�!~�Ci�P��Jvc�Rˮ��#� ���	b8h�⏀�[b���Fr<�18U�:3�j����������᭵��^/�q�d,���8�B��*%��&��m�_�Wۢ-Zψ_�q���y}�H4� �s	��-��mG�i�Cn�ҵ��Hv�0*�"q���=�� �̠�S&��;�. 3a�I,���x6"Ge�]��C�>��#���*n=�����L�ăY�[�fs�gQ������$b"i2D�8�G�����x�	?b��7���[�4�i'��|�I<-?��]Jx�c��|�c�+�>M�_e�z��uP��ù܇����'_��x){K<�!f Z��ƕl/�ac�����6"d Ü�A[7�J$��X*���k���[�d\�*B��Gt�56D<*���S�G�����!��?C�f�$������� ������=�¦W2��	Eɯ����9Ja�A�.�]�R0���ai�?�O�Hא;�:�+�U���\� �[��L{ޠ�O!�9
�7D�����x��袛^����n`��dsTf�1q��(���4��~$�B���ˮ���N��ݶZ��Hy�@�a�5R��p�pw]/��&� �� ]�W�5�`�0����v#��P���O��(aI�B+6F��9;MX��>��K����F����1��>/��"���Tv�v�=
ˣ��hޚ5�--rGX5u�c�{�A���޸ZCR��7G�8R��J*�/=�����I���j� � �S��<����ǛF�Q�5��߈$��% �ȭ0�F�r�}��
Jp�AÕ��d}�(Z^a����T��Cߕ3Ɇ{O�u�Vb9�r�c"�Ū�E%/��c%s�Y��C�q��MV@������&+a	��h� ���ެ�K�����p�}':Gn���C��&/?2�Z5_��͍����M�y�_��1��7 g�Y���~��h<�%����b]��F�8��ۮ�SN	P��,����&�^Os7�����]~��-�Ƒ��H�)��cg��& ��	�=�r"�����$J���4����)?!�y:V�!�W��ܨ蕪�+7n#�@L;���Iʃ�3���}'�{��ho3&>�B�7����b'�w�������niC6�^l!�!��O|���:�.5 3�ؽ-+5"�8 Q�Tj���?pHM�_���&D���I���a���uSD:�%C���6��j��TB:�6C%�o���C-��s�����y"υӪ��í�G���E�b�kq+P!4�>��e��.�L|�ɟ%�)��x�W���l�ν*Y�}�0��<�Hh�����#	�����ã��q��'��c����st��7N�u�v-:�04(z��������#s[u,��9-�@d�{�xf�X/_M6�	�i��1N1����F!��d���Z��I�2�j��M��_�.�r�sw�eG������)~ ������]x �-�y��:���`}�x*�.��7y�A�w����k�o#!�C0	�l��.F{NJ�75��b�\NX�vmy)a�4���r̸��ap����7���e�ڐEZOM�|a5����	����wМ�j"�Y�U�r�ﾳ.���'�����WT�j
�q~&������ȫu���O�H"��O��>Ɓ�Y|�rt�	�aGV�A�~s�e�h��4�|�lu��ܸ�i��y�M��#��?I9�$�����L�Ez���R5}�����s��dh��E��mPƃ�,N���e�kRi��p�Ksc���J q�a���gۗv�:�-����"Ñ:k����G7-�->0�r.���t�p�)!�{qo��6�J�pN�[��U�Z����� LӘf/Q0��԰�L�W���n1ĭ�1rR�� AȇQt�Fc�����d��t��i�Ha����8�!�
�<��D�-D��䴗Q��'E��?��6��|��'�)zIM�1�	"�&\Y�s@AJ��E�A6��@���]l^R{����Z��'K��f�����d�u�?�Lȿ!f^�I���7�6cY4d�0N�9����1��֜�R`�H�259�Ӭ��MHu����=�$H��Q�؀_rn�?c�n��Q]��<��L�tx�e��&Q�RMz�&��c��#K.�R_�&�=>���W�S�-Du��;�s��.ط�	
�A"�"`��?���'�m����!�s�����a��Y�(ќ&/bs4y4��o��G�Q�
�~�F٭������wiԱQ*H�/�2ap�,�'�-п�E��rswm������*Ԁ�"~Iz�EXǚ)蓚�����=����,}���G�C���2���-���lٙ�g$�ca�:���&��xE/�9���o�R^�x���Ą��E����#�m��Ӟ{"�;!Z`!h�>��YcY���G.ͤ+5$��5X��y�,���C���ƹp����0��p��pp�I2{��_���#�#;fn<�2���\����'��q'�8��M��曷x�@��8��aZۖ5	}��&f�F��͚e��jm�d�j`<6��`��-Z(3��S�]�*=�p�Ď
��4,`�S>e�y fu�^k��iGB��&?���m�������W��Iː�u]J��u�|k/Dv��&{�+=�yȴB����\��ܮ~�$�#��>��`��gƩ"!��3�i擤�Uf2���RM�ց�>�(KJL[��Ps�'�k)D���	���铚�h��l��m�D�z��d��p��8��ϡ@�C�2#"��7��ٵ�o��Z�9RD�p�H}'.�P�/c��v&*�\�Eǩ+c����.�]8Tդ���s����|
�褕<N�I�:q�ؗ�k�z������$6��p��3��iΈ-��_����J�JpM�!n�O$Z{������7�����c���%p�Eh,���`��qgK�Sjh@�@�������n����dQ��#���7�o���k�$!1�H��5��%"�)��Y���Sq�-�.�-C��M��~�I==�@>�Ԉ�[˸^V����QG�0O�F��r�7�� z���t:�;g�a,[5�x�I!я	@5<w�x�5�PՍ���"2S�6�#���Ȏn��<��\�ߊ�|�����̌lbx��>!�^���p�>�2�	<9+%���pz�.�A�� g�r�E�޺�G����5���+/oΡ����26�%��3X ���JS�`z,!)��4M4�6Z|�R,�+V=`GI!�Ӡ%���N��H�a��/Y���wB���9a^�Oq���f*����ُT0�l4I�Y#�{�����<����]���6��ԡ�0b=YɈ�|
	��)��Ԝ�jG������Y�c��5�����H�� �V�M��l���`a0�{͙D����+/�m��cDbWE��ǁ���c8�~�1ȯ�9��P���"@D����d
Ȗ�P5�F5 �A:UHW�O�@�\��.n���:�*�Г��rJ�#���`,@z���G�3���_ܭ��A�����c}��P ��f$Ԇ��4o���p+#ƣ��{�y4�b�E�_��TI��V5f�lz�6U�/ݞ���Y<���o��حcz�S�wy���\�\z��d t�T�ePf�Dc�|��Z���T�1���=z�� g�"7>E+/+6|�X��n�B����Ո��m�:���b�.��6��Ն��j�f-�"�s�>g�*�Y�[-	"�u�g�a�`*�H���p��V�T���`wr�q|^w����P>�(��'�ھx�n8�)-7A����O��ch�k����>�/j%pz���_N'�h��=�K���B��>�<H�VLo�癥6�dY#ǂ�S�;7;�7}tܑ/SmPK�*8`es�g�id�Cݢ���FT���-�l�� �O��I�1>eU!	�f��SSд�6��Һ����E�y��z��%*�χ20u$a�ʝ��U�-�}���;f�4ȯ�,C�>9jM� s�b;&P��Ĉ�)b�06d~$�MT$�N��'�,;���C�̼e�i2�E�ϻmO��zw?/��X`0I	G����)�7�9��@�W"��yq�=L�e��Cw{n�f�ԡ,f7���@����P�����X�~�Sk�`�0@����>S����I�{�.�*oF��5c���8�h���|붗�!��ot�;�!�&F���O~��j�BC��YPbt/wk����b�Ÿ
�tw��Y�+�p�խh�D���im0%�	����W�l$V�\I�+���%�d�
�6=mHW-�$h0��w����n��z~=l�oݾ�v�{���K�r\�<^]���#���W�$���&�
T��Q�D��4����Ԙ�jsVA��*�TG��@�I��t*�z��Cސ}1<�3��gˬ�FA%���� `-`�,w)�=��*����d*g5ߝ#O�r瘥�x�A�2W&x�3P��~�(�	����|��)[�zn���G�Za��zG(pr��Ja��Hc�l�>jEp��F���1-�mO4Fx�#"Iѵޱ�s[��9hi��͔��=�,���\��~j��IS�����gM4��#|���_=	f�W+��<�߱KAb�n�}n��
��-�Ġ&]�0�j5��O������J�<�QH�?ʓ�jS�V'��/\ԁu�/�HplIiK\ኒ��^�mj]���\1�n��|�S9ja��	����>]�g�,���߽/��D
m֥xKk�m>���K�shן���М<�FD������HvQ��K5KĚ?)�vx�l� ��y~r�?S9��b�Wd�x���;G�L�HJc>X��F�Q~^1ѷ�B��F���5��ħW����#�����Mt�2���0LlpQ��y�ƻٜC�:�T۫���^ßBup.ζM�	'�TB��D���o,.ml9�a�,lY���>�Ƒ��ב���	��vf��k����ߨ�j�PI�G���7���᡿�	I����у"�RH}�0�h4�U�R�%�@B�H���l�W�r$q���'�����Ly�
����7m��E�L���(.���,������b�-b����6�%g��	�Fg�����=�A�v��~·�,����݋�="]�%;x�?7%M�h�*r�n�����'�rɋ�X�o��P��%�/ζt���&%���ɤ�U������S��
%��u
x)?߇�-؃�$ʗT�H`����i�P�Y`&�O�@H��Hbo":J?�g� �eb�N@:�T9�]�m�9�|$�E2�IF���҇�.U����x���j(o���Z�H�P��WNܶ��{\��zb��KO_�|��͝(�cܵvMP�q�%�i��f�ͪp"�����'�Iz�����My"�ޞ~�u��PS�r���Xp%�iCÖ��-��:�8fJ�qu�d�y #(��u�Em�]�t�7p�g*1R��9{m`51��o���<��xN= �UV���ߍ0Y9/��mzk0Sh��S��?㧁 HU|AD�����h��я�D����b�V���+�@�ɝ�<9���+���b-��E(U9oM����I"PQRiQ=�7�+���UĹSn��z�r'p	/Ӆ���ܑŚ�H�,�|0U\�`B��=dA:���^@�jÓ�����K�<)�:���Z�h�9��\���:(��lO�<`)��Lo�mfJ��Ԏ�h�z�M}4��y�A$����օU��;�u��{�uJ���W��ǧy*vͩ�fA�|xȆ���22X 2V����!)ސ���4[c02��� �6Xw����MV=��3�G��������CY�Iwxz}:�{|L�b�U����yM� �ùkv��ve|�#[��<",��^\M�G�z���K�=��C�3��m)Q�ޢ���[�`cg#��DCHڥ��5	�V��FN�;h� � ����SǮ�K�()�g�Pg�4{~y7��r�}�2jt,����(����J|�����U	挈��+s{�eqN�i�dN���f�N�ƐB���N<�Mѧ�pI�5��WA�r߻L����e���k�P~n���_�	[X!���#9�f5�ܥ��
O�c�k�G~;�̖\�82��ί��	��0˧�g�<
�E�������nZM�!��ۼ��ӼX�cʼwU�F~kfu��$�~�6�Y���Lt4m�$��W�
j��e`�A��և:8����T8�Y]/Q6-s�_��ZP��]�r$��9�o*A[�ol���]�{ U/w��<�������],4]�݅ {{�#�[�'ݻ~�dc�{>gd�3L���c��]]]�ןUB����%��t'K�0l�>���������}yڪ��ڀt���^��V�!6�A�d�Fs���K?�cS�̤�V�b?�0�59
C�����q�wE�M��������u�\:��V��	F�*�e#*��l���[F�3QhM��=ވ����p#<eO�0-����+����K�/���3�7@5ew�x�����9E�=29N��=*��e�o���	�h����U��7�֨L�W�. Wb���ܮ�'�X��pDu���$��r���<+-.Yb�3X�ӑ�W�� Ƣ��1��
H�}�.c����`��:uΜL�T��H��1�Z��{�	.h.��@�����N�s$Z��uSiB�el����"�@�F��W�Ҭ�b#r��Lh�76���cj��%�O��I ����6�ŷ�ϵ%�4"J?M~I�U=�0w��A�o2A{S�zq��A
����O�hR��� ����a���%Jsja�/�o�8D�W��Mv���v,L����ݶ���cUg^�{8�I��U��2��d(��W��?���u���5=���\2,D�;���#�|5�l�!�r��]PB�����y5��R� >c=v;ѭ\Γ%% �������27����������L�����S$�?,g���(؂Q<��hU[�pd�P�� P���(w�s�o�j|t��AM�L�c���΋�������|�k�O[@�h���^�Po'='ۋ���1��n���蜧<�XPe��T���PI�wW����%��C�~Dm����JƇҧ��vHUN]]><{�U������+|H=���}�E�5R󎳝@�
JT�N~wR��F����g��cr��q�o�}/���7�ȇjXѓ��L����3�,I���˓�$V9H}	ٹ�.��F:V����	���=���|����ŷʀ�;���uL�ZS7�#�IR�a+NL-�$
Ip��L�W����y]X&�%����e��`�g��
)	��cs�/��p�{�~��|k9A� �Եh���V�e���Z�}d)�W�Ϲ�� ��O��0�-ǒ����]1�p�uۙ�ﻤG¥��سq=QN�L�m6t�6��A3���k�n����q��1�^�6
wc�:f��y��ho��j�1F���_\+g/D�p���/4�����T�.ϙ�P�Iôi�n��,����K`��C�A��pa���$�B:��Bw�c��M��Y�A���Su��k#�q���Z�c�{90�f�����;��a9$8M,9�M䢊WcC�x�I�SA�wHH�kٺ5� �um�h�ۚS��2� ���6#=�Ģ�ǿa?X3pE��l�˝,+��H��$g�o�1���Q!��Y�%�R�[�1)U߀]��1����S�f�`ZR�?5*����[�2�տ�$I�؀�R�eY&��̋���#kZ��[�o�|�`x���Se&�ѹ���Y���>A@N�ߜ��F������kE�]�淶i����V���e C=�m�'^"���N"��·��cZ���n\QA��=/ursbj#w�?��]���C'����\Ⴭ�!��G��/̏ܯx?���һ���HQF���{+|�6�ώ��	v����K��Y0����!̓��k��d��ݻ"m�6,?����]�'�N8	*`�5Em	p�Qܾ��t��XC�H�ؚbZ���n�@"?h��V�O���;E)�jX�-ٙ��FZ} \pg�j���/w���J���Sf&iUA��7� M	�g�dg�c��& ~ޗ��PE�?���7z�M`���^�IL�CE]%@aQ��4�#�V�M��] ù�^�_qO�8��g�#̵	�}"�b��@I<����u
6Tb#2���4c�4�J����z^�]����
}8ij��x�E����Xf �4����p��rR��3-٤���Ǐ`�JИ�ig�Ug�zE�L�3�UBYpX?w\w�B-S�@��=�i�u�MJ�N��	i2�9�K^�ګ����	�%�	��~`��O& fhp�F����~/U#{�1�b�kv�ԭa�����p���Dw),����(�=;�ŪP:VF��,���=s����k �:Ռ��[a� #oj���}�Q��@'�ZAk��o���md�� ��|���� =�
,R�����F��-�)%�t��{�dϣ=g��'p���o�M�\�'������S��oS-�8F��䈰$�Y�\��7�l�Ngʍ�$L�H�sΗ�s��`��I�O$���1���_~���Y��n�3ЃyV�^;�\O�)O���3`�6AǺ�;x�T6Š=w.�X<��ɵad������h!�BhD\�ʅ�� ��1Hk1f��}u~�*xbшz��_=���3F�&Mӊ�{�PH���=��=������~>+��'�V,�a��������w���x��iw�<tu�jC4z�h�J�e��T�Q�tR�OzGʡ⵨E�.�DAz<#[f�h���z�%�K��g�<�3G���IpBcEF�Ȱ�fGlOJ$'���Woe���l�%��'��s�,��̄b�U�Y�����]û��G�M$�����WM�Y��?$���x[���̽��y�꓈��z����Uh��r@�C�3
�� ��qϷ&a�3xH�!&��Ӯ��qC�TjmJu��QRD�.Z�ߴa2a�-Z�b��1�OX�q��	*�8���B�H5��R9��jeDQ�@�X1[��؀��h�.�l��x��D���:4����3v&?xcp-��;��j�m)I��)"|%�ص�Ԡ@1H�M��oq?W���/�7B߽ɔ�i��m	�
E	&�DT�e�0q�.+�T�U�a�3æ�׹��|�'�X��0�G��)���)�_�BÅ�M�ȫ@B�B���I�Q�_�v�w��	��A�YԼ���X�@�w\{9�1XIF��|2� ���B��6�0��b���܎O�ha���q$���ߡ�ż9��˸I��%�#ϕڗ&H�8�y��'B�aV�Ԫ"��6FO̫�BD{���_�>�'�mJ�%fs���Nȗ��Gd��l�zҚ��9��$�7��U(�j"H��J�}C�r�������F��qY�W��j�r���l|=J���M}-p�U�KӤB}p�O����D1��d~�V4S
�h�ьԮ��@�=)�@aOԬs^U���Lc���\-2��*~�����΍�=����jQ�I�S�Qy��͎����z��j�M��#�����+�|I����ԫhP-~�J5`��b��{�,.Tg�ߟ��N{������2�r�Z4�jX�K�����r�3�Au~۾���D��gg`���M���+�L]Q �U��Z̊!i��vQ�2��(3��hB(��lJC5�EE���S�G��A�`d��E�ʕT����}M�X�c�ez�S������+/���:!�b�jc��"�a���5R})h�2�H+Μʵ k�
�{�J|2A�r�{Hp�D[�:L/G"^�����zU~ű�P��C�"�<�.=B E�l6��G�	�X�]�z��z޶1=��zֵ���
r۲�eV�ɐ��'r�|�/��uV�πf��i��[�r-)-رء4����D`�2�	'ȳV��$*d�i�m�k��g�(7q9�׹�}ocQI��M��؀p�������v���$�U�\�����g@{�86�eߠ�3�-��j�:ܕJ�D}�//�����l�3T�wˡ��e�R�_�˖��G�N���u4���O��I��]���[�+��(MO���n�Є�������%��"8�t�|4�A��ƖL�M�=��M�	 �Uݘ���R�����yrPk�	�������u����� �k�R`�8W�0P4��Jv���(�ǋ��� ( :!��Fv3���|�ݫ�i���"�ҦQc�7�oнAi��6��I�Q�$��@�6B����0�����7�4���_�j��Zb'2A|�����Ћ�_��s�O�*٪�3������Z���4����w�ng
��a�����oG���T��3�x3;����ؕ�J���1�*+�<��'Q���:���
Ji����pW|Q��~E�����=}c86sGɋ!E}t[��u���<
:�Ƙ����}»O^�?��Y�����C��?>i���T��
D�[����r�?W�����7��!���0�$��۬�7y�|�X�Sq��������A��T[�h�I6F�ƀ�]�$���XWGC���<B�3Jp��+�tM�>�����/����]�n�Q�0�6Jf�)
�m��@%E�[z= ���+�E�B���X8w��E~9cʤ9T���h��,���A�d_�*�G'���T�)�]7��������_�W�A���H��� |ǀ7���#Xܺ�NZ��3�����\6��kjR\����jtdø%h��ܮM��>��o
Dɿ{s%����j]�aj��㙙�Z��D?�7h�]r�r�_���!6� 	�F�يYxoB�b�3ܙ�5� o��` 
5���V֖i �_P����j�������eh?!�#IjU�]���=#��&���6<�#�'b�������'��4 Nj�'Zg�(w��U�;�[� b�4*��b�3^~���r�
TW9��/-?��Hd�`�U�X�b�H�FO��������G��%,����U�o�D��ܱM��6���gҪy5�7�.l|���{܈Di�{��`f%����z��c{�>%A��B��?��B���
i5*�1�N��1��ߖ��L�(Qg�>D��g����b
>$��Y�i;:M�붶)N��mE�bN���g(�S(�	��^.�C�S�X���8�����
A�0��Nܿ�j�m�����p$��S����CN��T&�'<�"a�O���:��\�.����OR���W,�@�PCH�'�0��g������#���1���U8�*/ã3���{yj�k�g�\����`!uD;��dn�[C&�N��0��k�/�^�?�M��+�n��m�d;m���`��F���{�*���X�D��Ga�V1�L+;�m����c�AaE<�L�2�8���N�G釽�{_Y�� ��ߟ�h��NG��ƚV]9�ވi�c���N��<檸
�	����K>��.�YV��;k�*u	SW]B���чΞ1�ӳ��l�ۮ�+Bu�)S��$�qi8��Օ�+o�j�ʿ�K���<�X�l�+����>�(֢x��#J���^��W���ѾylT�����uiT�Sa��}V��O�1x��ϕc�isc�cn����|��A�P4�MˮA�9@���~��e���f#)<���*V���'�g��X�_1w�ni򀼄�F�zQ���^.��޼�:8��NՐ���Ya�~�]|�`�p[S�%�J�Fx+��܇�M��)5�OI0�x�<��O.�9�Z�	6�2��ߑ�[��u�n'av�9�*�b��ۿ\Ev�dN�>
�Dֶ��&��?�7�z����̸h�W=o�����a�:����U��ѝ�6�����C��OX)���$j�����8�%I�`1�>�\�s�I�I�è��ij��$U��Zj��&�PՓ�.�v蕤�,\�j
����#?�ױ>�v�	2$m~����冋���>|e��r+� Dj�<�Q��j�:N���
��=뭰E�����;�W����1��K���4na�.V�K�����՟C�v����k�,=Y�>1^X�`h?�Pz�4wJ���:��jP��暡e���
������'�ud1�1L
��%����,a���,j����E�D��a{��,�S�6Bp%��c� ����|C��Gb��%��c?&�S�p���b1B�꛼q�<�>�]�k�;/f�;>H��$V˨����C��R�������{zr���V���Z�^�� �3���O����Sɜ�=�2���S@Q�uOjJ���b18�Rm���e,�{������8U`s��FV��V��݌N\ik�;����EM�c�n��	H�J0��>��<[[���q�ed,,����I�<�OU.��Їzˠ�(��-b�;��o!��c������L��1�0i����r��8���9'X�7X
�
o�fPha_I���E����u�x31��o^��H5s�/�e�L�N$�Λh���xR��kP�s[�>W9�2UՋiU�Kx�E������JǼO��������c 	�c'C�������7�@�@t��>����2��ء���Ka���L>3Bz���\A�j��lk{3`�S�­�X�-~(*Lڬ˥h�����_��L��"��R��ƥ[����m��y��uQ��2R��t�b��F��鲒K�7�{8���Wv��f�-%ǯ^{<sg�U-~	�C-r辺�_!7q"�4~?�6��}
��S�3[T��5p�|�(�_�v���j�N��"]Mpq�O�u $��*���s?CuVs�j���DV{���p�(Ї&,f�#E�C�eQ{8��Ou�p�q���}�mQ;YQi�#����(���afT%�)�De9��5%p���<����KO��ϗ�Z�K\쭼oBc�g�
^�%AL^��t�Y�s����ޭ��
��UlՖi(��f,8qyѤŀ͏7å��01ߍY��,%>���k��B�Ԗ���aW��<�ʸ>��7㲝(W�UHoK��ia+��Um!<�V�`���N������@K��oh�k��ec���Q�g��ݵ_X?״�� _���?��+S2�'�է����Jn���h�tz�a�aT�탑�ĥ�a�ʣ,n�U�ѩ��-x���=1�d٨ߔ�AuCg���Z�;rT(�g\���ZB6 ���7��$`�,N�f� �؞]�E-|o��N��Q�uA��0>%j�s�XF~��q@Jҭ��lL�7#G�Ƌ�#.� pvN�y]�iڹLScJj�Dj�8$�M����T�o���\�;0���K�2�� 2>&�vZ��,7iCk�GE�ɤ���ͅ��?�N�սe]�M�e�lv��
.DZ���_���O
ͤ�>t�h.vT⥚�5{ߥ������r�ya5�1�f�f֩vbZ6��loV�պ�K�+Y���r�B|��W�zf�l��Y=x�֢ч��ƽ�~�J	�Q��7��P�|~�Yg ��)��OP�wK\�*l	z̺�{�(��� r>���%k��@˧��~_������qKϑY��.pp>��_�v�}{mb�J�x�P^|6��2oy�1W�V]|�BD$����R# �;����B��me�������j��d ��(�2���d� |4�ƭ��ނ v��w��	�u�K�]�2���&�|A|�>�F�p��6���vg��{�aB���,r�����p5�qa��t�;|��j�+hp7��/X�ٮ�h�Aå��q�cݠ���ޙ:8%�7,P,+.pݣ�fˋ�g(%���y��50�����t�X�yk%}��+�x�S�'�"a��}f�՟�gA� �++iR���#��@[�t�Ͼ\�&���iL|��_:wh~�A�`��Q{V�ʊ��u��7�|b�:X�������4xgh�L��A��_|_�T� ^��+>��o7���_�Ww����V�a�a�+��+�>g��M���9�'�d�r���C�<^`��d���(<z?��؉� "k�Q���G�����:P5�F2�δ�i��;"��Ü��*��K Y�⏢��X����� G��(H�O�E��
��a�t�-sa~�ol¸��|������N&������]FR�ǋB�_�t�:��	�e�J3͊8�ame/m�ًh�Ъ��k�H&� @ם޵/���s"1�ޟx���Q���i�N�ɣ�YD*�������Yo�tw9uu��l>S�3>R����37#�66|�4n ]:,�J�:Q����ѧ�/�c,���X��ͺ/�x}���(��;?�|��1�s�YqӋ��Tʞ7kI�h82�>�^�Q�N�`7��$�|̀�|=6}���pK���D	%]xEǈ��;�;�H�B�VSC#u�8�����<2��ܑ%eB����bh���5�F^�X�5yfj�S*���*��&>H����{;������*���4>�)ǻÒ� �jJ3�OyT}vy�-`,��JK$�c�r�d����9?���9��4/�0*{2�A��N�K����������l�qB��:�p�o�/5(��TTE���~��9�����U�u����I�����"7P���7��O,���km�u8��ڳtvS�ױ�����T�Л�!U��X�5/d���u̲�-��,>o���,��N��v�&t�G�lK:��.�(�U?�Q҅��͛��$I#N
�D��쬓#�����5�ԙ5�ãy��8	7DL~����!�S�"ȵ��3rc��?�*���%�h�L�7��ђ���>��@�>M���"y�Cv�/�R�UNg�t{T�Wc���@��a������6u�D�o����p��vx��=o�O���g���i5���鱣5�i�oЮs�Y�z?N_� n���G��� �{��9���g<T���L���W�*E��I-���H_OG�Up1�O�s������l�ٮ׭ �J[���x�Q�Ael�k��Z��v��A�2�C�ݟ�Jw���-~	�mQJ��[��V�U �3����An���cr7鱭<o�"!k�</�ے�ȷM$�(U�<��4DP7b��	�I�<�br=?�}&;���w"���d4��h���n�#�S�>xp�G�ݕ�(�֏J�f{��
��v5�Xc���ޚX���4c��ָ��wԒgȨ�U>��F�a��jy�P�}�c������r�8�G�;���n�#v �S���DLƼk;�]5�p8m�uP�/�E���~�m��+W6��$L/���>%a^�f���j���/z'~k� o|�����[���%/�e"�i���$�I]�n��pu�7%�E � �XǕ8�s6����=����Λ�h�P�ĭ��3L8��/���ЌĀd}+y��[3"W�U��.=�u�h��$Qm�n@�qy��j|�H�������~~����K��	���U jT�4�v��~˪\j�(��?18��|O�AǌRw�hd��Gcfp�ˠ!/���TeBH�+�s��s`���k�Ł �m»W(s4݊kiAu��RW��t}�,��ӱ�hЯr�
gӹ(Pr��{#l;Ow�>���,�ι zV؁�odd�O�L7nS��ͅ_7���t3ٙ\�2g]"^k�+�i⺻�iGG>����Nc�O�@�c���?�44W�[��h�Y;r�ҝ[H!��H���*�������O�]�vϊ����,�k���+����T\[�F��*aq	�Z��C���x�O�+,3��X��{o)�ՙLU�=?R�`�\��[s?�֕�,㊡��
��
���X����yP=xɟ?�<�]sD����2�	A\�(Z-�xD�dn_W�`�^����ᜇYC��5~�!1�m�rnI(�oR�������
#\�����9#:��e��A`9lHX���dY�`(nƗ�順6�I�A�Fn�>tb���@�+����G�~B�*=du�lVa���̃T=�,���0��9���=����@��:\�����7��B�,@1d�l����E��N�5 �����@3t6�W{q�P|��`<��l��h�¾��ƛ�6ߚ�He�[54�n_�[��z��1:�݈��"���[��h��+>*,$���d�lIV�>&�8!�����e�LSq�4���X�Hw)\��`�#�TE!���UU�=X����%W؛ޏ��)k���@��s?��$`ZvN,�R���*��V�zY\��X�oՆiTud�h�p��>1�t��$��ѐ�!�ᨕ���P�	��F#s���X mb۰�@)�|1(ܑ�r��Q�����.z"��$3�w(�{Ϊx�e+�t|�bM
,mq�2+,bU�wXNbj���.���֮�l�.)��O�h�BD�}�>B�~h�g�o���O��Ucȁ��'�fE��Y7N�Ϝ����u�%8���S;�՘�k��o�F<��l���m�%������K�'�ѹ�5�@�{6)����! ���x��U
�m[o����^HJ�Oߟ{�hE��p	� �:�#{�j���)�� �6b���n9���~���ߺ��>��PR�RDB`3����+�N<��bӌ�����h��S����nk�!�͸��s�k�<.S��z�z���6�Z�T+I=isKZ_$���s�?�k��2�7�o�.�T�T�$E
�'·ʣ�Y%�DH�Đ"��jLJ7u�A�O�4��Lq��4D��h*0�l�E�@F�ǹ���K~]o�D2���z�J��� ����/�!Ik8L�' �����|s�Za�dB����̱|��5FH|C�� _x�7�Ɵ�d.Dx�H����Y��/F�P%׷�	DX�����Ճ[<Z�J��C�iě��s�d� }h (�^JY���x��>oz#h���I���-�ȑ<l	���M�{l�ϋЅ�C����O�aM;.�,7Z�B_c��̚a���
�	6D�R����ӥ,߉Ȍ�}��(�H� W2o'yhXYRj��	eP�Ga9��t,�g��j�UH����W�����d�w�����̿��FZSV�wݔ ��
�'���Z��m��Ncw�m�p1`&�8�Q���?�+7[A�6�9��d����3�x9�Fp5NYy�]��!�?8�\���bP���>����$R����̴A8��nz�#�%C
�0d\�-�"ZL�,v/�9���ɧ�"��m��C��>�o��$p��cK�A�Q�h�j`Zk�8BR8��k�%��	n�^=϶\�$�[�p�^�Y��Y���g汿��
�s�b�Z�с"��E㔸p
o3��`´헦���L+~(�ȏ���P���50Qŵ������X�)�������i�s��k!e����I�0��Q��Ӫ$����k���}K��,)`��R�q�hY�����*{�ґψQ�o�޻%������n��X_��ߪ�Z�÷OX?�R��5-���H�**_�}ލ�D��&y��e]������ho@���`j�ut�O���������h�ẻ�	�*�uW���t��B3T�i=�٣����iԾ��/�R8��¾A�If9xp%5$m� ��z��RͺSڍ����C� �ѣqu�=�{
21q�c�x��?�9�Jڹ�&?���\� ]U�fK0h�n�8��95�0�]*�U�B��v�Fb��,4�����cP��qs�}c2��Q��8�f=2�H�~�)�B꫒�A�����0XX�zN��(���� �S�{�[x���fz���9��㭩|�t���τ�!���5c������L�p8�I`[(�;�״7�B��x��׶��$�p���z9���sȶ:�O�p�@^kj)UϼI�/�ǳ��V"��\b��R{��[}֨{�P�R+�����4h��1Ԯ/����Cik$���ЯF��`�v��8�/�0;�əO�M�12�eJp�CO���>�����'��O�HM� Y��D�[M���Q�G�BJ��!���! K3��ho��^��2���bGx?�Y���`�&�Տ���9Vf��r)V�lߛ���64�|߯0傡&�����k�g�T/&<�P�J'��V�gX�Fٛ��Zf�1��[C���w ;�? �9��<�V����xΰ^��s���=֠��>����=-��D�ݸQ:�;w��k=�B�y�9� 7T�bz�zxe�NؿM9�ϖ#"���2�YU�����9Լ�ϳ+ ���l�C��IS�s��76h8o�z`]]������_��,*UzQ�瞚�$W{* 0�����Q.of�ԁ�t�h_��g�4�⣨+�v5�����͆لG�SZD�k噄��*_�ӉVD��t�?���[�A)Dz|��/�[�@����!&�{�_o���v+�j���(�wSw����c��%�ݦ��@����غ���6�G�-M�jc��+��{����ȑ;_�s1�B ۮ����*�һxT�FV\���Zۓ�H3ڠ��T/����%�7R��{y4�V��|
��B�ӢŬ����]vq�3�ѡ�s��&��XH�&O�+�`ŏ���P"��%e�U�6���4�|� k�{'g�f2�ƨ=�fVlc�<�C̋8T����$��m#JX��̰�����C��s�
!~8���CH@�-~�Pv�q�y�C�`����-�Q�+Uh�6�ޒ^�s��;��4����T��
���v��c���)�F��K�{z���/���bd�yz���\���4�p���E֙,�v�rk���� ��(�GFLkR���L+�����_r����?��mn��wПNɋ�iH@���
�Gv ��;��S%�U`���!�uH}2��ȷZ�zy-+���L��ɱb:�>�R9�?������t��{��2��@�@�LQ3V�� ��oI��J�z��ٷq�cT6/���a6�	�/-X>'��z��o�kv��5a=cTN2�c�lR1��s�:;�����-��5��GJ8�z�D/�:�wؽr� ι���?�I����%�^��{�x�dA��v4x?���ok�,�* b����Ǥ�Ĝ%p_i���&P�_U���:�.�[p�Os3̂�A�6S��K�Y�z��,�؎R��*������|�n��_��6�J���r2ѹ���lI�T�~B����룎ћr��q��9�џ��T��F8o�lѧ�-�dr�z'��U�d�X��2q��%�l�i7���������IL�<�:1TL��{):�5	sfxK��7�
�a(BTJ/����k." U����Ts��GI6�%1���k(`���j�5m�r�]ٳYɯwqli��o��~Ä}�
{��$w_X��Jb�������Q�%s������(ԛ҇aGGz��� ��-�#
�"����I\w��+��!�����ZO�;�nF�{��fG�L}t"�=^U"}D�㚫�,y�ʂ��Z����V.�e������[�	4V�z'6%�,��_�h�f\Bj�|VQ�MQoD���D�Z&���4���� ��� ���a�ڎ2����.uU�����W>f�)M� S׍�7��oK�W����r��(�7ح�)vTd����0r ���#�H��0��B�qB@[Z�ڍ����R��E睃4���h������U���"�q�^ao���ּ�I�"a_e��L{�"�N	hU�[��r����% �ad�&��6)q]�������嬟bO��$��2�����k2�8�K4�E���Ȅ�H�#�:A:�!g�nߡ���!�ƴ%K�Zg:4������U��D��{�[�l���%��2�����
7�ٔP�^J����k1ۤfr��R�֫�� �?��hjfvHI���"s�	�j9~�Y�Z��Yr�?\��&G��\H�iH)�ӐhU��I8��6B��LC&�#w�87���=]J��ؤ$��J��w&�������m�b5�s�����aC+Og������G���`�j��ْ)����N�vS؉����
�Lؾ>mXr�)�dy0�%�i1P�ca���2���ʖF�N�c4.t0���I󘥍\hD�Gv��>��.���~ָ�oCa���T�V1�v��~7R	[�� �Q *W�M�nncP����z��ק|!�T��"���!f�Ss�0��ϳ��v��ș�b1��YE����0of1)���sO1�.#A��&�A��3w�twU��R�<s�ݥ,���V=i��}�����ȼ79{ �}=��2&��]/����1����:�O=�� "�������!����[�r�EѺ���^�=�Be�78ȯo����B��e�@�N���zv�=���2"#Jy޳�͈	�0W|�%�h��'�q���&&>���Ja��1d�6��9b��4�y��Q>9BKB��7�AF�~��q%ls�`2灙��)[�"{0��"As.H��|�pd/�݅�zO�$9֖l��pg�Vf�y3�o�y�-���\ta���1�x:�]�o-	Wd�Y:�,2����2@;p�AH�t�Q�t�CN+.��r���ȿq���m8�S��� ��w�5�Y`�(Hr��e��4r����5�h��H�f��	
f4��
� ��,�����8C�_}�k���J�kA�ɩ��hL�Ov��c����L�s��-&�ۊ��-���ųP���do�R$�
5^9Ӝ�aU�Mf�{�C�
��.{���j5�h����U��dK��U@�����t%�yK�\O7ah��;�_�/����Ol<�6�=+em�aGXl8l�2����՛����r�8-���y;�gb�����]ᐅK�j*��a��H��Uފ������[й���f�7rdn���.��j�\(�ƥ���FZD)�-WIb�����M��y�8nfV����({\$�ȭ��GE�����.Q�4#���7Вa]
`YC1�~���]�A��Y��7�q11���-[��l���A�]4�â1�"��0�kݠʗ���Q�z�	�]v��3�q�&	�%&<��P����"�ۆ�%�E�S�i�`�εC�T(�>}Ƕ`���,3~��^������#WϋŞ�Ֆ�U�$�('����v������u\��5������ϙ.�V`�+�°��oz�̫%s�B�2�z2(���2��JW^�" �&���'�ж�G��$���rډѽ��w�Oh��>��q�vQa�;^���	[���:L,H��l�ڋ��"�?6�hgZԕ��h�
Aɵ48�i�[����C �)T���7�C�#-W|�q��/НX���a,���w��\�u ����@֒����N��.�.�����R���<�R��l+5�rC���j#Lc��җĊ3l�C�$�4��x{x=��6k�b�_�rA�t27�$��.�d���d���z�W`�M0����}?�n&e/Dm�Z$U%,�9tWv��!]M��D���q��Ce���2�o2Y��Ig�hq�M�ʫ�ױܒ؆fTh��>��uE���S8�R�-ᕈ�haJz���@���Uʿ�vc��R<�#�kϕH����N<M�	�K"��JE��[e�U�͙��D;TTC���zeĳ�:���ns�'��.~�X@j����؅m�F�H���=���d�?�]�	W���/_G��-�T/*�"�jׇ(f(�}���|%��zD�F&��	��<��R
���op��f
�%��	�k\��WJ�3{t�/<g~}��V���)&������P�:���,mhn�ϭCM,n��B���؉ΨE��Ό|L5��1�9\E��v�*��,o%uI�����i����l����$�?-(U2[4#�-����y�9�6��D�d��0�,�������D�0�8M�=��?iL���t���V��Ӭ��]_��S�m��dKm~�.��պ��F���'��;�S�]h�=�Ꮊu��Օfp+�>h.B���=R���eN�+i1�"*ʁWt���J��j�IP�a_�:�-�k-nB��)�ΈN�=�������ߖ(.��E��~
�4d�盔��."���nM%T��$"F�]1O���mO�t֙c��9o�v`�-4Cc(1��;0�+̓&4�Ks�S��Y��Č������ ��	�d��d������dI��4��&
I�?��kю�*I
��a�YQ�Q5�$
ۛq�GGD��Ylg��PBP�t6p�B�Z�#�����[Ց��0�ޫb� �׹S��n�������K��R���)�+o��R_Vm1k�D���L�Q��p���f�Zw�h�����9!�d�L�fǌ|�l􈺦�����-�kG����*�v�ذí���P�m���!(ͽ�[�cB��({'�m��F�l/���%���S]M��� �;�KH�*e��y��`R=.X��U�q�x'KRBD�H�[\n{ơ����aB;��+�|c�C�)l��8r�-y9��UC��O�����e�v�nR�q�N�T)��F��M�MB�Z������,S,C�
U!�;����=ϊ�IǫҽDw�$��c:��՗�$"�	����s�s����P��84GI��f�F����]�lZ0����|�!oOU��n�A���7stw��mYx�7��&N5ohvM����dy�;��h"�w}8�i��i�[6e�8|�XQ�p����>:��������B��˛�iբ}oVF�*���9�¬�`5��_���/�8%��KV4��zכ�[
m�<L��r�MM�mky\~�\�U���*^ َd���U� R�zӘ"c�-��x�tS�9ƍ�O插�W�Jx�ne�TU��=^�Exn7�v폃=Y���y������hG��7�-CR�KP�8���q5h1�6r���εL���3zOIY{�ML�l��*�<0�'�*��ȱ�AWX<L>�aH�h~�
߽zd6�7��>t\�O�+>ڪ8G��##�l�����~5���G=��QuD��ӓ��q�ނ���\��mk@�æ����A�
5��WȈ�I�����$�o���@�C�����D��j.��_��u|Ls�1{Һ5m1���_�>k��N�a�V�����H���vڞ�6�\,PO���?�3>w�r5���S�9�.�� �L@10�����v��&�t���]�r�}��@�31+�d�hh�=A�C��:+�u@�P  e@��o� ��1��x�L����.FJ &,s�m�+���p�<`�ZC7�F56��mޚ�I�*�â�"�v����$z�N#��Ґ#@	-@�ڶN�j���J줼�60���y�B^���Sb\BZ��8��'�ڒ)�<8x�=&��k�Z��"���3+���>���8��(�_e(�(��In�s/,�DB�Y���̑zC�rtB�����
D�{ۻ!ϧٴ�?(4Z�~��Fu��v'�M���[�[!��k�� �J?�������8(MR�@T?:�e�J*/&<}g�YZ�(��{cƨ"H�'^����5�F��x�>�{&�P\�鷤b�lOƷ��V��R���C%�D�!S�����HXạʔ��b�������_�m�i�y~�ң���=R�Y>B��,ݷ���}�+�[��B�&~�=s*��=���	�C�0�v��ԦE���U�1�_��v�^�,i�"=���5�����O
y�?{Fa��o�l����r'@O�׫����1��4{��2+��I��8&@")�s���ھ��htF��̫�n���o �ҥg��e[0���4�vA�W['8̋=�p�a�RMZI6��i1qv ;$C P;�
����_����f�����b.-l�����/w��V}��
H��\��Ӱ�@�����(�W�	�o۠մ7_�Y�$=/����#�8awɀ�|m��A�o�0��]�;Fqg%��f1AP.�0y��|gm��d�_pv�>$ �Y��d�C�J!��%��]��Nz7k�An;�$�T�����ĸ�.�5�0������h�?�� ��?Q��yp�����U�榥�쐽	-PT
b���Q��N�V��Q��]�~B��3�[��	�6bC>��m�뮬~oB]�� ��~�a1@H�1} �I�itǢ�����b*u���21��6I}�Py����.�3�UD�g>��Q@>A�h��ݳ=9�,����j�����!Qh�L�M�@��^�p
�����&��Q�!�����T�aC.ړ�Rz�gO���ʵ�!"?
,���C˓dѾR�LKlY�1X���6Ä��Tۋk�!�~�'���NS|1��?	�ȿ��^i�>��}��ͣ��A�f����4���SNڤ��)b9�|��K�d�+�]��СV��N���9���z`����M9RC�޼�ri;�a4�Ydņ�Raۿ{j�p��(�38��UgES����E��%=śW�.,�W�HČ�5g�{k�*q�������mnNK��� {K��-[��F)�F�#���Qle��/���ym�.�
�M��F���t�5.�O��+h�}M��P�c">йĄ��s*S_�+�`1�Z$���j��P1�t��^9��݉N3���^T�:��gms	���������ѽ|Y<��cfx�?|��C3��4(��HJ���h���syV�kʕ��\�=��_�<�,7��H�W, �Qnyiq��s���] �	x��Uβ�����3ixށ�� 嵉L��
S��в�v/k ܣ��>��%�
�5�ݭ�����ǧ���k�Z���CD1d>���`�!�Ŷ&X�)NoBb5�&G��k� ՜H��t;�1�Q�u��Do�%"W���,�@^��ϰԵ	��4�蚶eO��?!���)�XY����a�tCE ���I��I����3�y�E�U�ޯjf��%OĈqt����kS��(�o�v-��-�/�Q�������Q�_
�o�~I�NcR�˛�d ,�)��\�~uay��Ơ`R\����d������hQ��df�)�u5��u�r������K�U���C��Ǎ`���T��9�X�[�W�>U�{���o�����J��줣�N1/��BϢ���Nw3oy����ǰ��zMoT���e���uS���M�C>�ٞ�4=J����͋�b41c&b@z�n��/zQjt����c��f?N�����"�FZWJ�7!K�y�Ӵ
 ���e ���_z����\����Q+3l\X��w'�(5�*��Eɻ+���,9��3� �1�|9�fӦ$���⯚ŋ�)��r;A�υW�F��^qJ�$S��m����\��\[!�w@��?�8�C�1@�Fh"���'M�$ϓ�O��
6"{���]��V6�+":�dd�M���"_u���Cԧ�&�Y���!q!�E/ʿa�Åh�T����KR��w3���^8��|���{����	�(��}�)rţs��,���C̝s�Qt{��u]��;������o�Þܮ���yN������"3��Z����4���W�}�Ea�uB�{1�ve�������}��@m�j|Bb��Ѹ3P���-��K~:������p�$��7$
��wk����զ_"���0�օx "�z�R� ����6����hI?�Ldv���/yEW嗅��O���j�{�ig�\P��g�t��C�x�� ���9���
�f��;'$*]_}����9�|�i{ �ε���.�<'��|4��j%�C�_��^W��58l���%6 ��O'��d4�� �O�"1WL}�-3�TM{�pxl��
_�4ȇ�=�L:�퐧��(�s�.P�?��NqL�=�F_*�R��^q�+a-��`7F�H���Z@%V��Ȧ�O����@���;�7�Eǭ�.�y�_r��uI��6&�"^�ԈY��-�U̗�D|��*��9A?ƻ{�:s������ѳ_�9ߕD�lB����L=��� �?�L�b©�ݷ��h����0����)�g������X��I��MK���1/���\@[�p���dx����&ܾ�p_�jY����+Q_eZ�
['�!�Q�\�|�O��n���C�1���q�C��	��C&Z��FA�iQ�tom~�w�v���Ɯ��9�#��<㢗��I�4�ϓ����!�W;@�������T ��ȭ�E>��T�?�ha�����6�B$.q����N�O3(K�}��6p�`��67q��RB?V'���08	{�<�/���B1wm�k&�b5�f� ;�����QCr��A�|ob��@�go˃���Us�Ε����䏍��������ȸg$��Fi�)66��������e���m��O�)m�}��̑�Jw���w�n��^F~]3A�G&]2�P6h�ښm�]�kb�߰��Դ�o!���"�1G0��e�++	��Oor�L��/�UP�%�B��z�����e/�܎څ \Ӻ)H�^�-L�������)s�>i/�����G���C�w�A���Z�t�������FL�{-m �����ն&Ͱ��+�L$G�Lc���1,u��``j1�2^�$��I���GN�����D����]t��in|9M�+����g5�T�oX脉ZRٵ�!�9�{~�8?�#�Ü�wiK'G�
��]�+�ja�!+S	��ND=�l9����1f�p:ɤ�BP]���	/��Dd��׶w���	w�r`o�%>\�"kS�������V:�g	��|�5�K#�g�(���Lh���Ufl������7�^�C�ݾVr0v��ȋH��� �r�y�o<��"a𸺼y���rފ��H<�u�s���CY���$����� :Q�&����y��$[��.�nN��	�b5�5<�f@�"Jv�Z�w�	B�^{�DsB[G��_�^�(���A�e�T�]"��1���7�ɡ1�T���Z�OK�}?/�{����&�g�3t1N������Akb5aL�E�M��y��ؿ�p{�lQ	I<�'*��J��GT���v'|ٍw�Dq��x��M����!�` ���[%��H��6���٢z%�'��1�Sy�ӧk����դ-`jR!�!#0@t���B��8��)*Y�9&F|�X�`�-���p�<�\���|8(|i��<#�n���*��3�v�0�c崬��"q��)�Y���a@��'	��ұ�RiVp�,��(��"eQ��q.7����� Kx���r=�u�jV�{����%hF�_Wh���-�K˿r��^�?bj��|������#&��k��,=��+��Դ��u�Ђ.���KcA$T� y�?�)�;��"��������!idčZAX�J�.��X,�+w&�h��q�,.O0�Xe�o3�O{e�C|Xjvņ=���"�� �jMݝ� ��8����f�)�r��!����yjգ�iE�G���"�ɋ�Z6W��Om!�b��9���2g��k\փ�ln�/Đg�M���d�?^\6yu�2p��D�.j ��_u���]t-_����r�n��GX;e#�c(t��ݷðuu�nR�-����GT|��Z:,w[m-���5{��'�`G���B�@ܙҡ;J#�˦��G�˹�4�L6�`���q���Z�Ƽ� �l��Xߟ�#C�{^�2q=��1����eX��W#W������i�ToI�9�F������#�b"��^�|��2�s��Ex�Tݴ��$���a�
Y���v?/A�Ɇg�֨vc8���N��.ff8|�w"�匧M�[�Ϟ�D6ڧ�|�ho	�s�^cN/��Z?R��,Iy�oVX�x8��mqIQ�E�%k̥��,[��9���u��`?#����bc���R�Lw�Q���R�~�j�H�KzhC7�àe�OɊ)*�C�r���`ֳry�E�_7m�ob^�	z�gU3��r�lAP(��k��>���+���v%�V�krŽ������[rS��(�͜l3n�6���̢%�g��I:�ǲs3Vr����lY�G�Y�ߙ.��Z��R0-���Yv$��N��tm%?UW�ӭ��c*ꪵ�|z�CXn~P�qI̚��n�����뿮?�%��{;˲*�W�2*=,�ٺ�<�gA�:}e`������g+�E��Ի��}�.�����d,����	����Q��t#f>�	@�w�-�:w<���M<@,F@s�FVu��jvl�a<� 
�����9��k�P���[���{����1��E-H8�2 /�H��?L��u���+�1�H��x��X�URxq�a50�F�n*��b���PQ���՟::hy<��<tZ���x�=��f�1�Q����Rc���oe�/Pj�_5/���l��8$��S&�:���>�&�O")�?ާ�����
>��:�_��J�9��;��$w�����U [�|��v��<ѫ��y���]�NHG��b��04�A����Cs����8������?h`lD�`/������TV�d�ī��@(q���Jz��w��xZ�����BtwlU��q�5߾��8c�@����$ }��m88��?�bգ��������y��Bì��x��G �uѣ+Tz�j9IN�qQ:g9ES4���mF��aov��Y ���t�X�m�Swa�p�E��{	�\�T|�wr#�i����n�-��n˅�sλ�Gۄ]�
f�δ=�>8�0~>y��n���^�x��9��Y�Y�GL�qź�֔�.�w�9$W~�*�8*\��/y$/"g;��6��`^���t���`��W��3��E������������)����$b�����`-B��Y�p0%׉�M�����{�cbic�8x�9 N��=��������bN���a	Jp���O;�	� ������|׃Q�8uD��\���ʑr�)a���z�[J��[{��h��R����+��:��䪸�=A��fF7�
T�J�I�
��#+�[$���Hӆ�"��	�K0��ΈA~s��:�SSyp!��[���F�,�D��}��mxs�Ǵj���M���V-�6��e+���Ͼ~�`�?�7� 	Q5���0�D>R1]<I%���m7��c�c�Оn���鞓2�op�\GY���<��[ â���FШq�]s�4���s}l�z�̴"��P��s#�U�3q���+R�O��6��Ɠ�+���5f���/9�*�����GW��	�4;e&�u�]�'$
����(��h҇M�{Ib�6��,OZ�����W�w��\QR9��|n^Z��^kp�D�����o�=e�P��JM��+�;��q�߼�}��x���,���(RO�W�=���=�{�3fl�Z�����%�c>9�M�^����k���n��6nrĘ�ѱ%�8wէ���D�W�knГ�B�#-)�;��H9�_�O�
T��t(���
��v�Zek�Ӎ�a�)��yC�/o6�����|l�e�z� {�\��G��R���b��\	ėr&+2��-rKl~5V�h�YV�������f��~��.?6V3"g>"����#S�I����~?��$e��~I�W4�`�Os��ȡ�^L���y��np��i��y�!x��,m��Y�ݲ޿X��[7D�� ��0�ϧ�u�y�,��1DiR��^��Ǹ����u;��&P�kM�.�n�����:���pkꜹY��/��{�J�w/��đ��?"��2r?��e��)<$���Q�M��9��|@�=�坻�c c���tXW�s8�n�"!���X�6L�pĢC@���<�J׫Ι��k�$��#�^�мq�vAπu��0I��#�F�B�瑛;�a���kV8�� ��̿HU���h�M4k�7�8P�0�u��n?�Y[+��T���KX�g��q�N�F��`|B�6�L^e��n�u�p��Ҧ�Hb���o=4�A@M�����sc^k۠�����Rk�mR/��ʑh�����[$p`���^e��E>�,��ǹ���(���R�۰��}<���+���P��X�L�bF�LY�O%��@*��I@d��N��� 8 �����\��H�v/����Cs��.�c'�+�3��<�A[�}���3��U�=��ʖxA�z��$�PD,"����Fw���K��E�~�Ƨ�f*{�Ss�Bj���=ǻ"��=$���V��dT�#�2�	����n�v&l�$n)�~:^ew'�TY�k�G �Ǹh��\Z@:0mW����%`ʪ����<
�?�͐b���i������HJ�+�T�t	8���i>�W��a���n@��/�3lP�� ��<���C�\A��0�p �O�1g3!}������]���r����� ���qc�v������O1�8�����#F?�G�ҷ��?�_8{��t�����ش�{���6�9d5X4 #&�y(6���I� ̧T¨v�GFD0��p�-f|��չ�|���URM��$,��'̽bﷃ~!�慤%�����L���1�(u�&o$]X$S�&N�z��3�Y�5��C��Z�[��� ,�e^,����v��k�s٧?+mv���Kv���u��Q�W��_���izuI��,��f�l�����=ĕ� �Et,�%���ٔU�
�ޛ��	
L�2�R�<n^���ol8y������Zp�u����S �{��ۜhU�F���|L��m�sX�P�=yE�u��_v�~H��6ݡ������~�OHws��=)�"��_~���*��gxk:�d�ғ>��^8i�R�Ef� >��Ǥ������#cP�୺y�x��ԵO��듲G�ܡB��p�x	?����ÞKk5�FWvZ���=qP�cG�2��y04�>�9���=����֢}m׏�6��UmU�d0-���Jt��k�7��!��x�7~A�	��H���������ZN��ks���~R���}�,�F��fm����Ė�wu>6��;jV�v��-䪘�"�h UG�mAĩ�dF�����{LC�D��+ ���HJ<��u���,e����/w��x�yS����� ���Ss~G�$!tYn'�
�G�2:BE�������x�Ve�J��J�Ŕ���^��}�4ȉ�&6		���X��ȱp7��`���bpE���x:f���8�fN�U�(�V&ػ"X�KīV�l�x�*^��ke; -9k;�����^�0�/ZT�"�qI�v��<�-D#b��o�����a!��&�]����	z�Չ���!ֽk��Q�8U8�}�z�Ȍ��f�#��cG��3u��Vٯy�$���õ���$9u��`B��.��2360D
xMX5�l��Dę�C/b��C��@Xlb� Q��V�!�.Eɢ�%�+k�w���3�oR�f�����O�^Y�f �lqǰ�a�'������No)G*z�t�� �5��¼��&;a���� O����%|��z�ۄ(߂[��H��g#�qE���˶����������o�O&T�� {
H�>sw��)�W:W�� ���2<^kh	�Zem�wȃV�c�� J)ؽn�9e}�xu�&�QTl�o�ʣ;6�`FU{�M��y�,rDH^���y�s�����.���.�O
`j�B�/��0/,�Q�7FJ5]�\s��� F	�f���PE�.�ҏ5A�WT�ǃ�A���IkXֲkF������}��}��ub�9Ku���H����{���ge��'��y�v��h�k�]6Z�y�F=t<؆d��{tiS8ÜZE��g�P�%*NCB'z�
 �9��-TO>}e�Ĥ�Mr��K�FQ���%�*��e��C�M�*��-�d��Q%x��%`�I��;��`��*`><�L����5�d���Ԛ����� ��WD�M�S'Z�6�繏�#TH�����	��:�.�fZ~&k^�|깫) ��v
fT1W2h�Dis<b����C������J'���	F�ĭz��)��a�����Ja/��h��h���Y�s��F{���x�(�v�Q��S_:n%�ˏ��m�ñmT��V��D�����:=��P����>԰}3 �G]+gC&B��Է8�愕�X�c��
Ñ���#L@RՀF�V�P���Gz�'��I�@rD��
\4�(m{�&���;ӠY��,�L�/~KE��\���`���;g�/�t�:�9�w�s��"q�G�~����m��r É��3�i�^��>G�y[���Q���N9���	 B�J�Qy��؁�4H��9��p��ݎ�cy}0J"�&1'F�}g��č�f�ǌ�)���c��q`��p{t�Qq��:?r��t�dL����[ٯj[l�J/i���pE7*4��r�����NwK��=����g�+�#�h��[��.���l�k�n<��3��Ѯ4���f�!+|4�,�
�!8A��x���1�i�b����X��v��&����R��D���������6XC����;�=�n�i�Ԇ����q>���p�B���ڶZ�f�}��n�I��1�`5'ݦ��g����o�qD(5(
���kT2f�Ǭ^%r"�F�|��<�����|($�� ѡF��JG9��7 �S���14�����༎X�Y��5�=0F�m'���Պ
y2���r��/�P����?�J���(\���Y�:¿5F[C��1&|pv�X��2����h9�z���x������#�>+���o���n�����C�?����G��Ɩ��Wf�/s�}�$�7��өU�5��r}֬�����? �!7��,�F�i:u��4��o��8�%��� ��+<)����3��/�<m�z�RCH�?VO�h�(��Y���D��M
�z��<�G�K��<��)\��"vZ�~ZD��F���ʻM?f�Ȥ��&�D��g�xqv��-&������"�����%�8�z�Є���S��"���j��&�u���\{���L̻W�a_K�{S�J��N���ν2��>�j�� #x<�Z'��>�=Ѯ�NYE�URh�q�$ۏ��:�w��N/�C0T�]��g>m�}��A3�X[5��h����  ;82+�`9�����O����Xo_�_�wu�<zU��"���9^��o%�K���_�BI��]
��!G]O�.r
�׶�d�ɑ��Y��L��ZU����v$4$�䃄��ExB���vv���j����0���œ���ԭ0��m`���r3��R)���@p��Xż��`�^i\�@�ɓR��X�d�ѧ��_\�=��Mà����H��1��G5X>���MD�"b-�{��n���)�RD�>nT�fJ^p�h*oˠT�����"#��u�_��ǰ�~jF�P�y����}��(� �=NB����V�Cf�N�J��k�Vm�_꾕T
9p��Ѳ;�����7��O�
�������&�4CÓ
�[W�u^Cep���P`��v&��+>� %�Q� >�%�c�G�*.��[8(P�p;��ĥ!�.q~�4L�fU598�����tf�Ź�q�����4����U�ɋ����\���˗�e��ʜS�n3�1I'������~Nu�:.,�vJ��t�M���;�f������`@�'��NwQa�HYǯl�9^�oZh�5XECy��S�&%.}M�ӈ������A�ܦ�"͚D�pYZ���\W�1�.c[e�0k���]&O�[�SŐ% �xo1Dl��'}ih7�Y^O�2v��-��T=�ƴ	���5!����01�o>߽}|u@�͢��󻐈�U�����H.ܺ�:@�j�\p.;�Ậ��p��A��Q���*��^)�����M/	�@8mHlf�3$��r�MJ�}3m<r�0�)��9���[�?��X����.�<��aC�dk�B��~�"�g�d%�R�i���� z��
��@��\ƙ������0ץ&"h������^Y�[ ��L�ɀ��JIq�AG�lE���Tی���hª�SX��u�:�l�%'�t�&l����q[�m����L�c��z̿���{�ڔ������df%��^��p��he?ښk�S "�ր��b�f҇Es~dd�>!T�9$��[J���g��_>�5ZKfɿ6�����b�!H���z��ql'a�bF�����mR��ܭ�<0L$אoxI\��Eg��:�*���J=�Z�l�h��y�����X�M7魀@��ɟ���?=JJ��[s�\�����v�jCܤ��%������y7�k�f�I��¼J�~���Sh!ä^�&�t_�]���HY7���o���x�>;�����&��ୖ��;�Q�N�>TJ�D����u_����,��">���J���#R����;J\/����k��%��U��_
WELf��冏���׋@Ă�W�.�0Vl��N���@���"�U�cc*F�=�˸ģ�Ǚt9�[$�ݲ����oɂɴ��X�:cc� � Wiy�M��[�Y� ��SB�!l/�c���L?zf�Ϸ�V�{�����ϴ�!K�����1�l��
�����|yx�(p8W�������mE�>�
[67ɿ�L$ J�V�-�͉ ��?��$1~�TkÈH��j���Ֆ�.`u�Ta.�l�g
�
���}���Zb[�~�u[6��F�]�]�Q')��a�CV��t��.R]~e#�ʇX���D�r���G�u�}����c �Iׂ��N[O�3`�j� D����g��m����Ȥ�+��S���<W���ID���?�ss�7Hs�Kp��$W�bQcp�Z�լSk����-5��?�M}s����1�����W�a�],�a��Sxk5\w2{r�"��(%�^��
���UX��\�\S{bj�c�n�Í�᥾$�!�e�a`1ag�4���fe�e9�!���c��ݭp�sP/'�m�����6�+�JTDJ�͍q0Ȭ�A�SZ�~��������ND)�NƯP�4�%���w�ڙ��U<������dt7�/�]d%6��W�V\�Xz�O�?5�>7�<#�YϚ<���U
��cۡ�q6�9�Q���&�3`�ί"ب���$��᭕� �30�T�3�y=��"�	-pݐ^8����u�߅�=�	�S�1�E>-��ء�?m�kl].����<���塄N�/�����R]�aV��YH�F�X5Oek��XV����L���'-s>�CF��p�'��E�����B��	����ʲ���&���k��,b�����Pk�t ����)`{�<!�(���k���w��!�nC��8��v����.�&��2�z]���,�XL,+Y,�Yg�P�@>��
eޓf���@�$��{�]f6�]�Nxd�iBٿ�K���{��,1�����A~X/b2X^ZV"���{SU>�� �]̏���[g�;"eu>�Tb�RN��B�g���u� ��~kLI.@m[������x��@�������$�gF�4, .O˕tu���?��ӫS��?{'�q��]h�*6�	;�S�W�T2��#v���n�>U��ʆU��-�̠�O�'�4K�}�{}�~���m����;��~�n������g��MJ��I)�k��{F⑀h����{��}�w�D�w�R�H�wVz��Rq�FA��g�	ݼ�Xx�4)i��	nT o�xb]z�F$-)�y�$mEh��Z�l�NA�PLd��Eĩ*&��VG�)���#��ߐiR�T�6^D���`L֒����r_�ybA`O�oC�n��΁�#�K2I��j�����B<P�T�'��vS��yu8�t��Ւo��~V��N$�J�N�2�0��-��Zؚ��n�E0����)�r+ğ��z۵�
���Y��3�q��=�:u�G?=���À^���r�	;_y�r}Y��W��txz�1<�~zl��vՔS��� �C����/C�D�7�i�2�pfxKP���7�>S����"#F�Ay%t���7�D��K�O�|��pR������xٓm[�o�y״h?a��P��i���˫�}OhJ�igj�J(��]QOP��ayk��*C�<�Ps�5PH����K�nYI���C�a��P��K��f�lx`��u��sd���Ӭ̗� �2�iA��p9cO��.O�K<�ٌ��D��ȵ�8��Gd�8U��l����	��\�z&�h�M��8���DMl��ޜh�/�f�"6���ƐK$����O��*3���$��F�Dnmoԕ)5�����.BrK�@k�Vp���vʉ)0���.݇�$���ݸ���i儿4bl�@�٩����8V@��S�Ț���L�0W�.��J\YJK������e�m��,N��Mn�wR�nq-̿2%f��C�N��u��լ�$��q���!-�o�C���yFZ�,�j��98��:ol�����ǎ@eQ�ʻ"�FJ��4��.��P���J�$!��U�f�l�%G+ƹ�ZAy:1��������ZVENJW�8����l��~7��)�@�%;d�ω�[W��\�<�f2���-�e�d*�P��J�6�D��������������y�����4b����	�&�H�4�y唘*)�9q�Ѱ`�����>���n��B�y�z�ݢ�U.���74�������V�=3@H����G��*�@s���� Zc^gD;��s���r�!��0���d����%����z	��}�kj�^_n�aX��x��v�#s��Ab�O"z@�Q���x�ڱs\x~�]IUB"��}�
�Zً�ݼS�gc�n��3� ��Q�3���s��%��J�a�7�j֠�w�PM�g�.R���&׿a��s�-�Ȗ�i����`	���)�Ϝ��щ9��zy#}Hg�)�w��Xj�:�b��D�Fi��^�.m���ɋZ��}����$�2>����R�yz\-.�=�*��Dl�^K�M}�����pw�����d?d��bj ��ǳ�+K @V	O|Op�/'������hQ�eg+[b�$��l2����i��|���hAj����'CM� J\y����2+���U� ������vZ�9Ҳcq�@~j����l�-��wSZPF?�Q���@�oNt��\+OM��^ʹ �$d���\YD1#J֥�N��]c�������tMZ �()��eW��{PeH)�*yPI*Z|�!=>j����&��a��\ȇ����:oc��	���wzb�H��l9��M��|�--�8�O�.����h�J^���q^�foPå^�v)ݪ�$n�ǰ�$�[	��^
L��G�k�	#?��iG򼓉X�ZsԖV\�'�%P���l��u�X.�� rX_�J��QTP����l����[���7}�Zp�0���� �|���w쬈���~S��X�Y]!��+z��.w�!po�*?<����y�R	4��]t��z���6C`����2bj�ᘛ�-�K�&h��I�⺹���6���f�6�������![��0���5Ip���2�� �_�c�j��Ax������h�����}}�X�oF�J��w8��������9��e�̉�aRȉ��O�[�aZș��Zf���L�vA��L5#,�@�@a�&e���Noہ�[�	,���.p�-̺�O��<0D�)������X�
�������nGn�p���(3���I!>�48�H2%�I�������q¤f�]{�摝�c�g��d�9�SA��d�4�yy�V�����BH䤢���FYVү��ũ�W�Va䢂��I9�?2�bW.��z��sr�Qg���Dc2w���1�]K�o�p<a`�`�?�{g��6(1L�IԋE c;���4�R���Eo��b��ЏF��c��:;��܂�u�+V���*Ԫ��������L^�$�L:��t���jE�qd/���.��9����H�\,
Q�^�NKHX'K��E럓�����3�C|����F; ̲��#�� ����1�*�2c�2��??f���&`|������f�& ��6B�y卖'����+z��YFߛO�=6�*���*�t��b��i��nd��.PE�����2�S���Ʌ.o�u�N)>y� A��@��z���X���V_�Rȏ�_Q]������|r*ܰ�ԄR�K�,5�f-���b��:zV&A9���0��N�U��	>w"@pK)��@"}�
����h �=Nm�@vs�sh������],S��>������?L�,��4T��3EX��Z,Wu<�Y��hǈ���)�c�G�+�nև!��IJ_���<����e��{�Ru�d��&�*��׀y(C�Iq�z�4�-��x�#{p9�E��<�j�"���n%�o��^h&l,-ݢh��J,-j�o_�,��-,�q-S=I!��W�X �J�E4��%'�հ��eC�u� �8�}+���ɧ�Өv<l�`JB��l��iz�WzASU��ir�ԋ�n?VR�e(<���X� ���U�53��u�V����>VY��1�Ӡ���3�+f��	���y�JT��o_f�é9	��t�7~���6y�C��jP� M��B�6��z�:8n�E��!¾�����Wf���Ү�n�p�a��8~�.`L������l�U9����&�8��X?Jʶ�8Ј`���
�L%b�_�ᜍi��10�(���c��c �Cg�|����X��m�~��qqQ:�	���%Zq��S�:���ۂ��
v�ӑ0�?��u���Ⱥf�s���yL�i|�=��M[����ܾ+fzy9o�N�$�u	��T����O}�$�O��-���qL�;6?�둰s�Pn��l��c:gt���U�^�t�\�D�aq�y�)ҧ2=/��!S��U%�iZq��O'��^6y�s�;Q���$��Z?pGc��˭k�T�ђg�L��i��y��2�ZJ&��ذ@r4a��C<�����і�n<W�r��H|e��iX�p��Wϡ����@�b�{'��2�w&2�����ɽڴ
����^�׺���1�kc��� ���{er0K�
���3�������ri�l�t�/���c|+���p�g&uq��2���
�� �Hf�'ᓣ�eIUC!���>ג�͇�����Ԝ�(���ǘKr�zR��>�_�M��~��G ��ZZJ�Z�P�����G�k6&C`R~>e����X�X!�J����K�+�0�SE�]l���tz��G�_��R�L`���ٻՄ��o`�|�q�*8%н�ؕ�n����\_�M�h�]�$:{�m������аQ��f�c�\�ꅐ�;�n�*�%�H�++�9q�'���
��NF��n7Ȉ7��7�|�:T̐
[|�5+�
�@\�.dS���w��4�	�AД��d�cDb=74�<��������I'�R�]xJ*�I��ia�+4�8�A����.,��5�i�:�(�c/��,d�S\N87U^�o���E+~��m��_&��U���Ѡ�&Y��h������{�-�d+�0���"
��k��\8��W!=���.����V7Y���y����'-���{=�[�{<�!d(������6�?�U�T����>����/&cÝv��m_7�?�,Jrs�p���5p��7n�]��O� A}'W;u��Ɛ���h�����]��� ��ID���m�ZL,V�}��.�a���y|!����h9���/]���� �%�A6�s:���x6��+LVɶ3�a�9�>ȃ�6����)�iblb��C!�{��?�"�sG��3�M���e��`��o��Ɓc͸%FTږDr�k��C5Wc�P�B��3�b3�M#���xM�D6X�%���� ��;�ͼe���(�8g6��wV7�M��b�����(X�焪�@�q���b|�UZ����%��3D�J�W3%����p;`+@/�x�b$��A�?��UZ����V� <�8��%,�#.[�����'��,�n�!뮑�4#%�?�Bu	�O%6�#�sV D}Z�$q!�q�A�\'U��l���N�^�Eܽ>.נ�y��ޮ�-�JYWE�hq��Sq�D�G�2�e=�H�=��ʕ�<�s���S�'���s�]�]�NG��7�ر5?���W�>��R��,Q�C�O6����_[^���DT�08W\Z�e@]1�T�ޛ�L�k�vi 	�W(�r�`N�z��Αl�c~�C�J�>vP@3d���jmx���8��
��&���@�ﭧ%��+s����1�,��`�Ŧ&�r��U�˪�S��cy���iݦ�Y6��/�<4��lN�(�)��R|&Һ�̱�#���H�N��!���f����f�A�Sa�N9N6 ��)�[r��kյ.�������un��B 2�k��׋�g�Ֆ���!W���J"�i�Q<|p�6����7�� ɣL*Uؖ-Lg�9&�#Y�����y���*��	�9����"/
�rR�~�gS�+�Q�Qdo��dע�S	���m�f�օ�~�uׁ�V&'�x�������m�*��z���bamiKo�u����1;��,O���Mܖ�W��ʼp�cٞ��"܊m�F�UeL��;����I�7e$ΟxbO`�����^��.�_G�M_5�&��@A���g��t���q�"�"Lɇa~t E�G�qs�\�,�Γ{��Y�K�>g���Y��!���?☕�#��qW����t����әn�Ⱥ)��O�}pd���@�f-ٛT�g̼����K�|���&��$��z�-M�h/'0�@�$�	(@0:��c�a��ӥ�l,����J�+q�z0g�֙�Cd��lr�~��_���a��蝀b7.S��$�i����tSk)n�9�:������'+6ZN���/����#{�i
�U(�X
E��<��Z1�;��s-z��[��*�ߔw1˒�[�M� �n�v��wP*��А'�j0�S��
3K��<�(M�U���ϟ�M�(�>����'3d�����;%F�;��l��}H7�u��?�9���ǵ�8ɏ/���i,1�ʰ�~7d�����\e��#�J|}@�9�Ǉ.I��Cwa�c�ڽH��4X`���Rs���}�B���`U�0��T��31�I�������]�-B�_�����g��D�W��&�r����6c�}l#��B��62`�(��f��V�s$yY����_t�(�v]�#�!���j��4����l�Rr��+<H��oE��NCE�aLv,ٕ����1���ʓ����>�K���l|8�3� �����:�����r�����)�Q'Q�+ܪ%��K���ܝw.1V����4?\Y��&���Y�|���1�"�S��ω���y܇�Az�Z��{a��:�w4`V�����RW��#���)f��كxerw��&��;�
C�u��VWP<x�}�~�0�v�}�aw�'3~�|�� -��Ϊ�:6�@>�����_Ux+_������}�\���H�oΚ�6�I�)��1xM�+������,?h�>bR������G�m�o�����S=�4,[	�,�{.��y�E���<����d	џ�4xC	�I"��&u`\�@�����mN3�7@Q�\e�1�)whN�wvH���w|�5�"��8J��I�|!�Ҥ��L�f��r�t�@�q(�a�����V��Pp�˿)3d�2�K���[��� ����DC�|��r�����}���,��;�/�K��x�LVQ������`���lf�`�0�㙇0��a7��=ª�v~�ބ�"��o�墐�!��~��3B��VU
UM�g>L�3�f���i��x]&I�g�����f���X1_S.�&�eb\ʅ��^��c���e�� �r2+�<��K?����?{KL������&iMw��hW�-'7}��c��_*NzO't�A�����K��ɛoƅ"����^���J�8�5���B���+D�H�L'��1=e��et�[Q�ᗀ��?}LR�����d�*�{�h�f�+*x�jڪ���7��K�y$<�v��v�B)8����ɜf����n�|� �D�ON��m���Ю��������[I�_ɦ�c�*d�]��b$�jl�&uR�M��@���,���0���ڨ7�&����p`��i�'	ޕ6�t}(?r<-��kVƫ��e}������6�8[��bK��}�T/���צ5���
+�:Jyd ��=��S�0m��V�Ӳm;S496z} ��3Mȸ�m�[aXy��T]R�J�f�TN�<w��k�5�Ne�{G���u�����4��z�]|�!�J4 �ѓ��0ŧӳ2JZW{�W���&=Dp����TO�����1�mB��{y�͍�+i�&�����G��U��&��(j���[+i����H�`q�
��̽����
��\1 �ڔFN
���΂/� ,����X3e2n�!k>Y�)�ouT�xX���ލZ'm}��c��1M�;���O�A��OB+Y��<��5��M'e��_�N��]
]�Ķ�h��d*�22mn�5�[g��.i"u��(m�q��z�'��!J�kzk��y"`H���8]DE���Eҵ�lp�ިĒ�]�F=�3���ز��G �gL�IX�$4w�u�x�N�]9�]�?L�Pم�mQ�;�T]Q��mu��;_��F|��oLz+>�*K
��P�@�Z�-�&F����$&"��nO���~Av5�:��Ct:%Z>R��H̈O4���G��\��q���P�н'�b��h��~�Kѥhr@�����՘�yc쯗	ڢ-��ORC2v@?���ã��&�J&���F������*	�tT�nN�.3#�O��T�QR��m��{t��&#=�SՊ�ޮ�Q��t4/k������b�cсUO��s�t2F�����5$~c��u�7���1���#7+�2N��m����~8%�C�(0I'�����P�'Q�P��%˰%T�I��I4�����Dw��oEe�Y�WeO�s����m���J�Y�7NJ~�y��lh�H�b���[�H,�"�ߍ�X��C�y����"[��M3���z0t�P��໪���w}r
!۹�`�.N8��[&-�5��8��淝 �A'��E�z]Z`$YSr�>��.?<G뚵�/9HH-^��	[�B���1�ݢ��nz�I���@�89tB.c�C�Tj����+�'�a���B5�ܠ�lUZ�QQ,LtNM���$�B_`��v��+��`Z,���-C��2��u��w�m�婤M����`��i�._�5t����$A��ܩ��%=���IZ1혍�J�n�O� �r3=���{&@HB�� (�DĭҴA\ך��Y���2�E���z%�*�8QQr^��D�$!E�QF��n�d�I�r�_`(�gl�Y���F��_����>lXV��E�>]բ���R�1`�6�P@���Aiꁥp�m�!~�@���M���6����D0���p%�:|��<��Ԝ�o�2��f|p��A[dX�����g�T�vm����Q���f=SB���Fc��V���䓴���E����\�:.���c�i���̥�g٪� �{%(��r'FDe'Uˠ���g����;�Hs틼K�[IB-hU�ͧUG��U��r �}|�;T3#����t�j���fya��gL
�x�8�~�tO;�Bȅ�Ê]ߠV���ȝYwZhf��
N�Y4�6�v�c�~^�Y^�u�'��~-Idb�$F�jY�0���(9S�)6H2�cG�Eh��^��@P�r��y��@`$2	}��c��!xZ��2�;i�^�+�D�j�W���ks���5�xȮ�)����]Rp
�PZ��H� UB�BP�V+���`b&(�����@M�zf��s�ץ�>����j�N�=��ޮ�����/���I(��~2*GE,Ԅ�X�ƕ�Hˮ���f�*>O�}�N<^��UƁd�F���o�V�Ev
��;l�w������k�ΐ<�Q�۵��bmJ/w�M7>|���.�������q�fw�V{X��M^rx5"�a4'����0�C	�h�x�	�/(�<�d�jh�/~#��,�ʶ�'H���;{f>��3+1j,����
���ϰ�ɕ�}*a#)�tŽ9F6�?|���iZ��#=*��R�^��
�5���gab�������p���k��a{�L�3:��1k���O	#7}��*����i�����o�qr��!OM�d�Z�.��I"�3�z��J�11Oy?j�.Cr������#�����8����<��!C��le>Р6�I�m�<)[|vYP�í#;)�U5<��j��9�mɰ���+�8倬,�k�)A_�� �ZZ��αUƣ�S��i*��
�W�4EX�J�����-�G����*�����m_�Ig�3���G�x'�c$���Rj���p����B4ʒ�q�@����*"s��$����6<�,��vAH�l)l;��To��|�������R ",r\Wu�c̀؏y��q�D� ��k,>l�p�������kl�Āb��)��a��w�C�˕>HWcd��/E9���[����҂r�eG��x�p�L4�a�ʕ�������V�7\�Z ι�j�^G(ǔ����R�{)0+K���P�*�L�9m*1�����*�c�a�-�Hl�.�17k����·u�]GC��,u���8{��ǳ��),�ō�P�i�w�W���y�f2|�VxD
�J 9�N�E
{&�l��b�=����3ЀĦǋ+Z�e��	�6��:�AӇDs��q��`��H�`�%G��EB���K� M�mj��T���}���-K�rpnۊ�S��x���I��
��\�!s�s�?��R�������y�sA���ʧ��S�/Z
������Z�ʐ8o������r-��^���~�k�L.�i�BA��:��.��Qq�k�!����04x)�=�B�N�C���d�(�3���XZ6�	�o�q�&�.�/��qE���Q��\�_r��$��X�:+�-�2cB�
���dȫ��k���n�S�D�z���PM_Y��>��rw��q��FN�w)��x���#�%��d�~��E] mq$����L�@�v4�uoc���l
�B��
�3�A��3���H�^�{��Qh��6�ֱ��͒�3zZa��!m�a��P��B��a�cr�����-���М�ղ
n]��)�>AZkB.]�0Ql�&�bCj\��[ c���ui9�=�?����[ ���+�qD
�L�r�z�uPDԯ�[�;�&���)5�(�`H��;ㅏ�"��,V�
�l�V��$H��������1���Q��e^96o/�]��yqQ@WF�Zc�hm�7����qa­��S��T��@�
�*��Za�d������X�^�����.QP���W��اA`1q��P9�|)ݓ,1����%�'�Q�����=ݓ��E �SLɝ�R��N;C�������e��j�\�mVPx��|�!~t�Oz~�*,�
��=#6�72��M��#~�k«LWle��t�ߢv\���̹S ߄�D���}���N���Ue����>��!Z1w�qX܋ռ��Q�RD1U�Y��%WSNm0Wt�{߳x`��H���/]9����/�C����f!�\�- �^&fb6cMob����RT��KoC4@�H+Q�s�'��S��.-���{#��x���hp��!�{\�V�(�Ҝ��X�̕s�a��_��w��w_55+��wfڇ.K�}i���u&�Z��K�Q�~�a�Ǧ�XI�%<��h���ާ�,'��6�'g�Ǩ�������u3��a/�/u�TU\���h!�����
1�Β�M�te�<g͈#jum����:���--�]7�]��p��q��;�ꍝFceF�ڀ�0���jz�|Y�2p��`_�!#1�Cڳit��M3(�{r�K����I��~ �[��M֞�ۆ����H��]m�A�E�}�볁K`�Z�+�����H+Ih_!ϜZ���F�seԤy
g훢�"ߒYk�����q��>q-.줕BH|i���؃WI�ދd���B1�:y�:a�p�`28�qS�z8}񢓣#�&�x׶p��EAo0�1W�������+1?�<�#�>qN(<��,?Z��YM�����)�&)�E�4l��%�g�#�" �rmz�Xu�H�N�����q����&���dz�T�F[�#;�Btpm^b��1���/O�c�vB\��6@١�|���M�nlg0��7�l��7�� �a}ABW�9�i��6�"�L#��['�RJ��2�tA��$^@	Y��մ%ڨ����r�iqB��M7#U󣓗H��#���1=����l���������1 ��{O$�ф,X[^c��j������M�K��V+��
f�J\c[D	�C�_��v.���C��D4��h�ȑ(��QX퇦5�zH5�S��N(߀�C!��;���O_O[�jDDƂ���J����R\�Cv�ʧMY%U�P��El >����!'9�P�g�J����wi�����5gA�!>P_E�u\�@��B�eȅ�ө]�2�sٳFW�$�4[*���#
�b�hʛ��69��r�3y�ec��,��W/��W^�ڱ&o�K�tJ>q�#��&Ɔ܀������Q�D9���Z5A������E�^Z���xz�zB��Kuƣv�]�GTQ,�ܝ�=�Lܺ>�,eo~R������ -�c@h#�k�
3��	0��!a)ë�{B�R�� [F�������
qSk��$�_î�&4���Z=%'Ank��Ćye�"T��ב�'#$^b��ɘN�1V��)x�&z�M�ŖE����ak��M
Z?�=<�M��Q�|Y���௽��C���z�5���� O�_�^H�>0� �]<Kج����] {bu��G�7X yd����<f�q�����B0
�׷��鷉w���^F��ze;Y*�U \/ʉ�DӚ�ۦ�B���C;q(�#0ik����\<vGA���&���j���~�1����ߚeX)Y\�]1Hl�`��.?����Jbe��wR��mw��,��-e۾������1�B�Ұ�&�L�N�u/���"�] �v�e�& �MF�ٜ�B��9l��`8�l�����K8�0#t4yw��]p��	����+�Цf�7��u?������S�e�=�NNwwf�+)���ܡ�A��_e'��C���
æ1���\gZ�������.�]�W\��V�=E�Eu\a��g�J�*���Y�(��� �^�h��;��.�S����GE���������'���UD�OЌD�xd7�����H�����=W�VLn���	�w�`����ɿ8*�|8s qY�d�/���nZ± �|��|p�}*jx( wm{c$R��7��MY�)�����q��g���˵�O@ۗ��p�yU��׭Mq�^; p�x�B'�-��=�󰵓o��,CH58㟂c��ӳ��[��O�K��[+�C��A�m�ʬ���&9$�V��E�W!jn���tҜYU�>���h�/THBF��Ռ���d@u�� 0|ڱ�(����I|(�&AX;�����K�H[�@�W�[�[8 U'tCG����k�b:�t�,��w�1��-��Ӊ9i�
�ϢG���߶ӈ�fL$a��~��wG�Y���Z$R����l�fߦsx��&���ȓ��lOv�����..<��+A-S�)}�@C�2���>����%�0��c���ӄ��ٵ�7F����ɽ�7���H�e~��,D"2qyͤ����E��f���Q�ecy	=Zo��V���I��~4YR���
��ވZ��P�%u*���2�l��2�$vU�ޕH�V�خ�i;�����Il3q��+��
�r�mʌ\��t�n���YE��6�W�?��/t�z��Q=L���g�#�95�ɵ�02G8��`�$�*����9�%6���
x|�T̛�C���pv��P���T\�lPz�l5+��׷���ts#����;��u]�ʅY�q1��c(�ɧ�o�_�m�3rh����6yf�Vu^��Q�{�e���f�����bj������)^���\�ed��cR�~V
�+�,uS�d��KB-"�WA�I���s��F%^�fDMA���U
��4�=O��v@KC!��d8�yN/^����C��WF�L3*�<{@K��^|@���F�[a a���K�1���bGO��7.%B��7+&5�X�pP��cF]Hl6��3R�gք�#�Υ(0���qk�]0�Um�	UpN%f�2��u'�Tc���o�V���,�2�/�F�m������VH?���Kǩ�Tw^K4���0�"M��4��B�<8���Β�L&�<�G��k
����g��kaZ���$԰Ur
ZT�^��H��N@c�1��E��{2cg�a�M
��0,���ޅ�ȦI�ƞ��Ķ�w�X�pTã�����nuk\��ֱ�41L�h���K�u�É�V"�8a�o����.d'�7J�{�|�땻�x����7/ K �W%�&>Oش��qc �L+�]U��w���a>���X����@�w�qV�?+56�[ϫ�I��ɠ�4L��* �tm�����ԋ-m/��"-a��NXt{`�<����s=�LUp�d
��%���PTz[�}nR���)���)�E��m�Wy�0&����X-^0�ɞ8�y�;�����s�ν����8�YVM6���Ԥ����f����F]��v��x�5RE\�0�g[�k�+	��3!1@0�9�l�I�9�0��0vlSS
�O=	TL%��d��8�4���j�lA8�
�2o�[���2 ��Wl#��b�2�%��&,�󐛲�H�Ň��k�J�w��\:z<5����wA�yZ�뮚�u_@{A�t�Td �da��o�mf���.B�����KÌ8�F Mq�!-�z����h�aR[��% f�g��y������c>[15���Ƀ��Ր@u�5Bdv�;��`�F���r�W��\ۅ�9��2�g>l���A��\߫$�
���{�q��+%��Т�[س��~I �8j�/�%M�Sjj�$�w���Ѳ�Fi��G�47c�#8����*[���F�~����}���;� ���F@#Fyٺ$���:�<�,9�G@`⼇�+l�z����]�YF'E��)�v�7����tlH±9����bSdu����B~Wh~��O4~`l����i�\�>�C�&r���׼Cv��N��̞���H<�@^ȗ�XX՘+�J�t�]W5I�wDx�4޳(CoY"'s)�kc��I���F~CK�<ّ 1�@\�ҺDkA�~𺌞�qØѶ��Yu�"[�r�Ya>��B�Rgx��~a/I�&���=�(ga���-'H��5�4��/.�dN��̴j��g�6���?K����/���q_�"��P����R��<,Ry���#?�Tcs>Q��Iҝ���o�@s\��#��wΣ�IM��n����F! ��{u wJ ����'���#C�<2.�k��r����^���HA��3[�iqD���|���.���3bW-YDn��C3�0u2U���f)S����'��U:�sտ@��6g>7����?I��u#�p�� S�l i觜ydz���Ge���<ޚ���d���_� �֜��^����*����~q�R�%�4�kw�{���$0?�,Q�+� ���0� ��o��K��?�eA�Ae�#�3�tg�B��EG`���q�Ew�m��x6�LQl�J�(.���c���������[������]EA5��0����r�4C��1��G�x]�dY{���K��hU�Q�6l��G�%�c����{����O�}r�j奇<���y���+D��ri���'���/	�'��P$w��R���T ��͙d��˴�jT&� ��)>�$o3U�U��;7M
�Ǻ��&��jG�:�Ӧ5l)��[���z���}�~��u���En��r��~��E���eqM�����g�X��0Z�oҩ�W۹�)w��GԻ'�CFG���W�p�"�N�7!�q*��oX�ׂjަ)��8�%w�n��Ysrkd� ��50m�Ew��jʃ+�W{�'��v��#���<Y5�u��8�z]f�w���V��9K�$��T$ˮ��,V�,��P'�'�l�6�s����̱T��.N ��6>b�-fܹJe��X�9k��5��<��Nu_$���Pu�mm�'�݅�Nm�K�����Ej}ۋ}b��fM�"B{$��XC~�>T�f7�����*�����f���E`�"�WKk<W23&��1�ii��~����g�7�q��;���pj�� ��y4� lG�{{�p1p�o+��{>S�R���L�@Ly���T���cQ���s����rR��:� v	�?��$�4i��T �I|���W7�����Fѩ��r�F��{���܎B�Z�e3vp���dр�zo4D߃qM�!�v���_L��Wh<�qu>��K7��)}5߭B.7���u�oT�}}�)��Z�7��z�f�G#�7���`R����ymt��V����C�L��;��^��o|���,&�N����N��z�^�1���f@ ���\�9qW�}W���`�1��Q��r��s�.��;਩���ϲ:������!6a
��' ����GS����P�U�����,@��gҷa���|�^��?}����/m��BG��
�~�kJW\i�߽��]JKA�6�.)��1v)$@@k�e�J��Ȟ'l�عa~L����Xܴ�7�������fOģ��#"?x��ud��W�xE�;-������o'.��(ʿ�cpPx�i>��FIvj)��7�aɼqwcX�h�b$�J��]@�0谚��t|t�U�=g�K~�g�O/_�g���6s4�����h�K0����q6p���mc�����en��yx�=��h��xcX��;A�������w+���h���'��X�����B�=��	�d�{��4�J�0��9�'*�~�`�E
?vu����MJ�}o[TI+�$Q���fV�w6��/̍ y��[o�Qv�3�7s4
��з���C Q:� ��24T��kwᅳ !���ð\o�֫�Zbg��Qq��M�4p�K�@���� �&�_{�HX��US铐@ )�У���}��:K,��7R5(�7�r��v�G-ݶ���t�r��t�t���6�����5����/g5:�jY8r�O��EB�;��/�\2�i���`U?{|�W��$bfS���<V�:���,׎Bq��
�R �Fաƀ��������	�=���U�I^�����`	Z�:[D~�xx�4s(��ۮ)�)��R����&��!Vg�����2+j$��`�S�߉�jQ�Ob�&� �t�a.�'��NWlg�OA+4߁2	1��;�#�8�����x�֝������)���@e��VK�!�!b� �nq�WE�!U�	뺰7a�Dm��#*�%��r����I8^���an���Bi$=a�9�>�� �MC�lS�ա�Ƒ0F&*���;���g;y_ڹ-�w��B	*X�XLsq�h��҅���U�ɵ}[�xmIc� ����vo�b�_��/����q�0
O ���D�������_�Ǟn0��5�%�0>��s~����s�Vt�-998g�3����/�5�KzM�
ե����m�-Y�xI������g�'Êh���QBM��Kl
q�Z�ok̏�1RYRLkW���I���$%oPz�h�o.7'�3�ML��F�D�
Fd�Z�W8]��EKV�����L�)~E K��j��Q�̸%p�~���|۽<�{ή���o@��&<\yn�JԄbB�����\S q�N�����R�Ɲ�,WG��4̌͝Kܡ���Ǚ�g��bn3Ǚ8U��t��.Y���0�b�XOl�+_���H-��� ����f��?8����gh��ÇtӱD��	����G%Y�mᛴ%���h(�F�j�P��N����c�ώ�t7_�*41J��#ؼ@0��a}��ǣ2Nx����N\LJY]��[Ύ-���,��z�$Q��M��H�uoX�6ik���}�!h�.T�������u���L��B���1�J!����y��;�y���c�V����b�J�.3!+���{�'ro'��#J��p���i���p6%�i����c�^˜j���$[%y���{�_b*Q���II��f�;����I�y]CrXnG;�F}�t+�� ��6�dߍ��tL_�K�R�!�0�$��O�?�W_�cTu��r�ٵȀ�>\����� ���s;������@T|�&j�J�%�En�d�)�)%SM�,�l5� �C78tL�熎>f{u.� ���H��4�t�J����bu���x�r;ƄIgz�g*^�y��#b4ǭ�ȳ�{�"s����X���W�xk�
����@����~���;����> ަ�w��?��!���bQ%����)� #mo�1M�/�Q�Xc��ȯ.��N	!���v%]wa���9�/6�_8��3�dK30Y'�#��z0�!m��\���Ɇ�8 �̊=���*��RFX�S������w��� �(%����Jcs�q���oI�J_��CpI�ӢP蠨�J��v-<���`�](eg`HOЃ�� �mP����x�BZ�#k�3 �%k���#�����y�g��\��}��K�{7:/m���ۮ�������,�65�i��&�őՂN��ިl���g��h�PK�o�*���B	��]) ☓�A���Zj���7��hk��ν����L�"k�}�c�o7I �z����:��k[d(�47VW^�qxn�^����5����BtB���c1!����]��w���֮�Q\R	��"�q \��̴�A���P�ա��-F�e,�W�=E� SZ��O��A�w�z�����_�U[A�	���Qw��}Z�ǡ�����/[��E�\�G�k��\�DNK����YG�����x�^Q��[V�v�EѶK��9c�Eؖ�_v� S�Ut��ec�k.��
��E�Տ�Gl\}m]<���T�ɰ]Zq@��)�� H����;�0��v�~wHR�y��EB�:�{^�\>_LY��7���*�^&�*K栈ؖp�"m��N�AKyE��K�Ь<���W�����h�S�@T��`��T�&\].��U����L������g�ɞ���W[3�i{#��J�%�鏔�]�z�Q�V�)N�R#�m�)�]�X��"3�;��uI���e�S)ƈ ��} �z�+�P����:'�72�[�P�[�q���^X��� ���o����A�R�Y7��Akϻ��f�����_$Xfn�b�xs��y�&��mxQ�o�XL$w���Vǔ�})�g�Xl�U <6�;�y{�7;�sjk�zGP�N�����:���L/���J�3�i�6�k���Д�6��R��my�s�q�G�8��Rg�)7�[��	�w�57��B>�]r�!�1�Hÿڿ�qW>�:"9���3�j����;��V�йA��LgG�"��s�1�u~gyG*D�I�]+��4B�w���ېum���-_#LM-�;�����,���i���{��TiN!� ����Օ��=ҍ[�"S���y� o͵g�U�^�:��D�쪃����9b�D�b�= �����ٞ�U�Kor�yt'�3
zz#��E�[�U��y�T����O���fuA;^f G�3���;Q��r�h��AML�xv���y����s�\���
R���qٕTu&H=�����h��o�t�f%m5��I���~���(&��桢@�W&l	�Pb�]���*���dW"`�]"e-�e���l��g,���2���R�VA~�m.n��#�p���Ɍ1���	C���8w�~�[�=�q��=O"Μ��t�π����%,�.�����@H����w�|E��(v>�ӟ�����2b�$�xB��|��dF0�<9��'�����5}�.���&�g{�a�Ht�Bg�r�,:c�B&���ӗ�_�HN`��aT�(:�&�H��+�Ų��ӯi̣�g�g����>�ck��Sg��'�8��x��9P`~]��}e��~�9�N5g������L����YKM�[wy�,�r�UCu^��lP��tV	��S��&Q=k�{�-L��{�%'}��"@LkA�e\�D���%�ů�b�ө��e�41�Ŝŝ��p��s������8lT��U%������ɚc<�ؠ	�Yn���TTд�����/c1Swg���"8MyC�o7Z5�F㷇A�t�Z�t��:��)"�'!�i,�P@
:�ق3�@6��7��ӞL�5�4�N�U��0u����G��R��
VI?l���>�#l����"���%A�#4�j{��q�Qx���aNBGlpt�8 P*�1v)D����������&{����EX�4f>"3� �_TE�N�
�M�ڏUV�M��";��b����h1w#�#�8�1r���{�wC����e���,o٤�I$�m�V�ʬ�^fP��>Ηw�o��0�7i���"�x�N埐p�	V��s�M*����-։ ٌ�� ��⢰OP�B;;5A�����6z/�q���R��
�U��[!(,D�[S=�Q	[QZNh`*����1��v �"��a%���7J�L��Oq�K�ڐ_Һΐ��R"Ŗ�g�#,T��w�)&��v�b���m�����Q�!;�d�[�to���G�����%�`�4�Z��f�r��RZ�7{�vw��g����u��$O��B���S[^��W���!���G$1]4�Aq�i�RU���v�:nч ����_�Q���y?
��ퟠ���M0ކy�[�K$���'�-vtcl-��22SG����k���YzX���U���Đ�}��S`��"3�;��,ᩲ��`K�Ҫ�xF�`�`��|�I��,���!��S���)���W�}>E�$�.tp3+��|�:����?�4�M�ү��Zfx�*��Le�\_���1:e)2_U'�Uhy.NX��`�o��:$5�L�s����9���)��NC�{��~��6�'5F��Ӯ������c.!�M�h�3�i�ˋ(N���г���!��$B��΃(��證|!1�I?������c9ml��ȱ�cHȢ��.�
��QRl�@���+H_5�����N���`�v���N���=$�J��@"i������`���:#'ْ�6/�X�C�.��
WB,��^t��9d�S����UK���\P�MI�2`�=�k}�A�5|�>���Y|�_b���]0f�`�"}�8	��l#�����rH��E�Y ��ސz�R�z7��d��AS
����N`�B|��/z��4?��o5��� ���Z�����C�X̀ ����U��S�9Ru�P�+!�qZ!�$8a�?\��B���
_mc歳z&t\�[=��9<��`�fo�e��]@��~}.�+� ��JJ1b��;�Di�Eew��o��:���9���P�+�>d��3�aA�M[">�=��G�U��'}78Z�Vo�R���6�>�^�����^o�zo}� Gߍ�vR*ufXide��N��w���t�Aw`J�@�˩����p��`3B8�B1L&U�b��*#d:T�&�{��9S�f5}�e���r�0��ցH*co���!:�K{:��E����@��:����wf-��:�q�U��A�^�������Q��Ml��R�R�QD�FE{��Y����u�Ǐ�5vS���:N�AV�s�^l�n�2��>�Wӫ�Lwt}�Q繮ZwX����wmz���Vx������JY,�P9A�@��=�H��k�${˦�NE�s+i����[P�$���Z�۱\nU!A����$+��{[�*�/�3����� �*��������#JJ^���$7�'%q��*૷��}.���O���B��_�-�_{��~��-}ۯU�'���m+mP��yepګ�!�⪴�j6��=���L�1��遥�	�~����أ��/YYP�W�s�K��f����:��k��������j�ԕ���#S�Y��{p��D�9v06�EB����ˍ�P��'=TS�1oo��,ҝ�ީ�ɋ]��:����Y� �PUx�d�Ð��-��E�xOIq��-(E��ë#=?�N;�)Ԇ�m�`zW�:N���}��:��K0��I\���@n���"�5�Sȗ���_�[)&�3R�D��X�-�r]Gma��]�w�:�d�t1�e� w7�C��MA�+T��N;GԻ���R71w�������|* �W�*w���;�r�*1V﹵� ME� �`ޘA��
�H��B���h5�uSk5�*I_���e�q�D�'�evS�.e�̉G�����@Bb�0~4^�;k�m��&�5_�c�FA�${��e���^a�G�7r���ӏ
���a��/�b�&�g�9Ë��$�.��������ޞ�M���
S2�X��2�p���6W3|��_N_��{pn
S�	[zp�����U�9�S�z��	�vg�7.����6�j����^ťc��$���E�ę]@$�A;Sz�À,��U��U�?K����ݣ�L"6_��7
�Xa`,�9��Ur�C%V�l;Χ�sr�E2���&+��w��"}����5������a���W��cR�{F='� ��_��hH֬����+x�U��������R���~�\�דa�_D��Z�CXKI3�A$F���_��=R�h�q\S$��x���4�w�h6|d�(��8wHx�J��l���ގ.�O��@9��h�Hؼ�F�BaH��v�Y.�2#N�{�0O�_Ȭ7��N�O���!8?̘7��6 ���i㽌+�lV]�"qt��7)	�zh�����H�
����ڇ�XK���	��pi��Ɨ����:���Y6&����d�( H�Sy'������>�� �Sb�w��P�T�s¿Z����N�ˈ��%^ߎ�9�)�����5�%±�Z�O/&��=E�t�5�Nw��'�	�zf�0���u�7��_@.��*���2����ć��e�!!�V��p��#��<�w`�kܷE�������eJbs�=b�pQV������C�8.⠄�2��=�67�^*7m?�j�xȉ=orqčE"��0P6��
�&	��2Lz�8uE�B��G��`Vɤ}���|���w7!)N�ԉ_ƫs$�**�z�u4��M�רV1�Qw����pn!�q���e�������(L[P���Yc����sU����K�<��Ǿ������0t�
��ؓ��/�f�g@M�ϒ�ɝ�#2PB��9V��˧�Y�+Rlb�='�	8���[e`8m��,"L��H�x-��̝r'ɵ`-�rL /��VTu�d���Q��co�����b�~��'�8�D6{qQRZW nEpC��.�����Q4�譳�C]?Z�M^������YǾ^��	s5v�o?�i�)�:�Ҍ骰wf�z��'oALg�z���g%3Pb�H***k�Ӄ� ��V{��RO���7􊊮.�-;W�� �;���
c���'�5Ru�a#(� "U�_�1���l�;s��䠿�͗!lY�`�����������eE�P81m�Y|�.�¶3���5�������e_�L���Ѷ�t�k',�J���c0ˤL��O,�8j�)���Q9�E��ru��$N��
��ה���9U��λT>���Gϩd��0�)��x7w2�4`��	ctRޥK��� �|�(d\Lpr%5W1���Ȅ�����4�u�x��6�q�N6]E������ޞE��B��P�e�ç8��NE:��M\:���[��%��aTl�17`������ƛ��0����q�-d�i ���=\����և�<��;�}#{xzD�)�!��Rt�n��8�3F�N�sU�ZC��8�d^��r����r��fo�h��3j�X��5}ކ�Q<�c\��B� !�W6ڷbH�F��q\�p^8@l�M3(#�P��8���X���
+!�_��)v�D3�)����C%ʉ!{.����r4�Aߝr�	�����z�`&0V�/}4��el�(M~0_�@.Y�����To���Á�
���m!���z���7!%8��9��f~�2��u(�p�
���P0���̉��X�]�[Us� ��"�%
&�C=����sP������<��4KR��<��y�7��vȍ�d�'3{����:1��F�S���dw
���dƴ���7I�*�I��-����	�o�q�&R��� O�)'���� �q�b?�5����ҍK:?����(�����NH��26�����
����Ev�|+��e�v�$w!�t~ռt��vM�H��@��UY��i��D�L3m�V���bz������r�h��]������g9:�zI��������=N����'t�1�A�(ǒ ]������OXv�
~i�-im��4j���Z�t�Eg1��$cW�X�ϝN�v��w%dt�W�r�|�1N*N��ՠ����	[$�Iw��7SɄ�����ܧi��U/�0��Vy��E�eL��`��,a�?Б���v��q�<v��r�BX���(��m���qX�Cw[����H	uci�x	U�k�6r��{E2�\�=�Et��;4�[�ul�յ�~5�8���lo�$9��f.�6���#-�#��8Jنw�DL	�6��Ib�SQ�G܉���P�٫eԔ�D�H�� �m�kY���lX��m�A�ok�L#M�i&�D, ��j��d��F#7g�3�y���"��^�Tr�s
G�����[�5`<br���^��l��^�T&4��{0@	����B�:�c����5m``���\�r�2U�����1p���HEh���)q	 aO��x��5t���6���	g� "���E���R�?W�~9�p��M�j�`�� �����)��>�\Q��,�21	�'�^�|{$�&�����$̽UG��x�|h�U�WM%�ź	8�b���Ar�XSa�2{�:��[�dt��?u������
�-_���9{'!5t�����SF�8ԓț{.�U�wgU$	 ԣ�����X)���_pJإ�㹗ƀ$+f��Ƽ��k&et>n�D�E��y���A���k��
K� _ra�`�+�b�Ֆ�
	N���NV��A��G�5W��=B�)����D����gآ#��	���s�	ȀXM��\�7e\J�����Н�ܩ*�ã�%3�XR�Iv���2�>�GƬ��)�pt�6�>�#����O�*i��5A�x���T�C��t*{��Z@0�;	��C��w��4
�<��zѲ���l��5h�_2~j�3f�ն�; ��$�[D�u�pۏ�Ɠ�p�r�g);ys�{Q�[C_�@���$����V�k�;�[�6��������[0܌��+R� �/��� I���	qj�@��&�О�K��K���w��y����v���*Q�{� �/-,d�)��4�����X�h��BOPV�>H\��n�^+?q7Mr�0l���X"^O���?��q�9�&)���e+�´XH IK.h�*\ٞ}�;�t�����R!��b�G��xk�?:�uD�^�v�Q��ـ��"�g��>K�6���}��yec�������b��Vg�� �
�FP*�|��D��K�j8�>�P���1�������=�+|�T����$��H��R��L;�$9�)�0.l]�����Ϲ��!���ǀ5 ���ߥ�q�ʑ���s��+w,/V���*u%=;�o� 6 㹜>T@l�/��K���V������#fG!�#�v�G��n %����t�����*�.�mջ���T5��������|���Jy�U=�l��4d hI���l/���)|H��st����y�JI�'����B�.�d�0��8���,� 	�Ó���!{���gW���7�� uϡ�jz�2��+X�^��ݟI�Ǎ��-R�����_�#�����Iָ7L8mG������%�Ę�M��a�U��
�W��ZWc���-�#�/���K�s��N���s)3�8�k����k���Y��,
ӡ'��ª�7Z6��0��W�R���]�To�i�����ͯ���p37���:�g��ϘH�2oF[�������� 6�gE��}B�2ڞ����y��"[�\s�1�Ȼ6Э�z�H0ɯ�=�P` W���tq��Z�%�	��ޜ���C���:�CD��e�ȹ8n>[�3���ƍ���S}�v�]Q�����"���SOV(yk�0m��F��H�Z�	�yF�%�bw���n4��hpe�/��dMU��o�'�\�,�Vq��F��4k�!�7��!�+��l�K�{6X��w��gy�)�O��7��1�������j�	kk��{����<M���݄�����_�%rEb&�n.�Fu �	����0{�-gHZdcA	`l	��Uw��,�g�9Uz�h�`)��I��8%$t�_�9ޑ4[ :�:�0�~>�Y����;J�D�d�9���Q�ʻ(�٨�����*��N5�r�>��1��S[Y`r�K�m�w��D�lJ�Q� �S���6��c8~����,�h�j^]��E.J�(��{l�x�U^���W:w�GPRPv��T]:�"8�T~���X590.p�0�c��3� ���I��T�у}fK��^D��C��qI����I��<������p�@��x���|�@��9���x�mT�y�/��b���vS�?֡�tSyHkr��Q�n���}<�S�G/]���ܔ�\�(LD�Tl�����ك:{%�\���J�D@̄�7=��8��F�������(��-�+���peV��9�-C(ag��BRd�i�Ͳ2A&��^U�����GN�Os�(r�ӧ�/�s�m�������}^�t�����o���8�Q�Z�/ݰ�f_e>4��O�6Ioc���v{��@���&��Ѡ"s���QN��9�Am�_D���u�h/����J�3�:=Jvp�:����r�����r��k`��:.k6g.�	w�^.�֓xme
s�=C��a�ly��$��#eͫ��]%zr�S��3�cr���ٴ~�dr��C� ����F�M0�B���H��1\fb��a�*��\���I���m��+�����j��1�qMc�)O�� ���b����g�0v��Oh�`Ӽr2��%Ip{��ZcJ��J�8��Ju<��=62+"i�^���E�av�$�{ctk(�ґ��R��Ш���@c.uE�'&)�w5�� �/����&����q�1
��Q�B������U�?Yw��0�*����*=��4�&2��-t�U����,�ⲅ�3����q���k_`�As
��)�O�-D���D��,�(S��F��H�ˠ�v@��m���E�NÙ�ԡ�[U刑���} ���$��W\�I$_;Q�Y��c�h���� z��p�0=���CA� k�C&xD�}�+ʓ���� ԣ�ǯ�s\���0ء�,�n�"i��@ #˾Hd;5�ي]�!�!��EEk�Fg�6^�֪�)1�W
�3���e����:{�O����>!����|lQ�d΅��{�C��)Ӌ���HN��P	˄S�$��,V�*�x�eѲ�r���tk��8'ծVW�bl��$�dM�	`��n.k2��g�J�]���c��m_��P�W��<�ܶGKdvwA�]�a8+da�~�kV�w�=�2O�U�fy����8���sDGf}�2ۯ�_>9Z#�p|�������!�Π�'�x�~��&FZCk{Y8���uB���
z}8�#._�"U�k��H0����9bu��^��+�|��F��,��d���-�\c\{�'�]��g���e�Na�B����5��Pk�
�v�����C��Vd� �̓)��\��>����!ISc{�M��J�V�Ic?���hh ;�,�l8f �G�	`�$��g��&�m���ƙՠ����c�R"�g�)ȫ*�b�SZˈf�gf*������yPd�
�m���ϯf�eQ�*��]�I��:�{^�௜D}���Z1N���f?{�/^Z����{�4E_qCh�^kl/ ����~1-P��d"Y����HBL�Ǎ��O;[¿Tљ�6U_��:�.�2�D-A�&epqTĺ�7o���+4�bhb��$���#��X�*�4b�#x+�I�K������uƒ��i�Cm\}${���_�Fv�w.��q"�|�0���ą�+�b.�@P����S{H8�r���r}@}'��[R�}�눙T_�_4��Q�G�?���~��Ȑ������:�%�&��Ĳk�j<�ҝ���-UfQ���@�Z�d�ݣE�2�(���E�43�d��^�WI�88S�Z����qE�d����ԦQݲ׏��ι��3�ur�$�gI�;����
6s�w��b̔�rӆ�K�0v�s��06�Q�$�U��uE_�κze &�1E1'�_�:��\y�}��`���=��� �+zx�XGA.�0	�0(�	��B9.9�U���af#�E�>`v���I�$"�j���+=%2���*h�a_���Rd��m�W��9'����g$ͽ�ڵ�=\�.�(ؿP�8&���Ab9�.W���~����D#�ǩ&����������c������sF��0����0�Iz��#(�Ő�{����[�pW����w����2u�9�B���1�e�����uK�m"�N|����F�L{���E�x-1S���4��C�-z��lQ�k7�8�-��zX�U삐������]a�ZHŲ��oV����._� _�[��W�F8�EM^P�L��3�{���Cm���&��F��QYS��6c̫��p���K8P@�hӕՂ�AaK����E�+�O�rL���8P�J"4��K�yx.[@T�l���"���5�	%�ۭBw�c�i�O�>ߗ����<{�w���d3��X��A�!��:�tLy cA钶�$3��j����Y���@��s�����?�q��j�(�,�#��K.!�G�v�-7�	��C$�Ƿ�^Wd�M�����Y�Yn1c��	�V <�ޝ ��W �w)��8���wj��SG��,�-�L�ʲ�i����YT"%�O� )28_S'���Zl��[,�I�n�d���=fH�l؝ ��ָ̡h������e�-lW��V�; �j଴�!@�0���X �Y��Ĭ	r�Yo.��@P�W�++�!Km��$5A��l	�w�Y�Y�8�rw��p�����K5�F$py~e:����;*��7�
Ϭ�@��o���UO�աE�],�!���1�%*iC��T�K˴$�A�ՅW;�X��_�?�KE�q��!2$_�x4�X;rg5 �_�F �'��^=%��ܴ�0X1���sNX([�L
ƥ�5rQ�Tr�Bȣb ����i��۳NJ�1���a��Bsg�ܸ�j�YSHvL��Y
���r�Q���MrQ�5e7D���w���Q�n����E�3^��� �XK1o� h1��T϶D�Y3�YF y��q�XG<h�h�<b�y���pQLL��2���D�SZ���3��4PjGn����rȳ'Lq(�qs��듭j�6����=�`���qm'qUOfG�WN["�  ��U^4&�;G_u��-��@���:b�U�zW�I�zU��$s���L�l�xb�v�[ƻ�A����rQPk��ACl���9��p-���%��C��%��1�!խ�����\Ñ! �R����M��ea�|S:��c�����͎�)\'�&���X�cJ;B���N9g�?�q:]k�a�#��5$J�&���}��G4,3<��Gl�d��r�=�7*��0�:�|���!MO�3������>(�~�͖�g�:r�Q��C�s�����#�b���>�l<��v�Qr�wD�[Z����U�g���6A���C�)��3!�#� ���7�bElvk�pz��z6�0���h�*Z�U��a*hlH�U���tD�A�Mu������'�h- g�~�RЂ��i�T��Y�c>{*� v��|'�>��B�����^H�3 ���ck��d`��X��^�[m\INՇ�l\��ڲ���478�M���C[Ϡ�ŴY��^0�C��"uzD}���4޶�ox����P��k���[k.�:���ޮ�&<�ȶg1������;��;]L{�������Y�K}�\g5���ۗ��cԼA#��Mt3�b=���r14�¨�a ���*�_:�A	��^���#�n�� �o��c�yRp��|iBu��n������2��h�d�d�(���P��x�W�̦�t��ābf1hE��-����и�fs����RF��Ccm�WQG����]��"��j:�`�,���4��py.O�I_�3������u�������=�ߟ�#��3��g�(0J*ᇜ8��x�P[LV��@�sw݌�Ո�N�n�-M���n+��JS6��y>E�h%��\Z4��c��fTE%�LN���\	���x��vYC���\d���\m��LTT!0Uj�m�ٽvb ��)\�c�	���łw8�l���]��@xU	o���(�D�K��C�n�`�w_<_'�|����.�O�ڪ�i�s�HJ��Q��s8��x^�u8�^������E���6���M���=�"��� ���ϿZ��n�-¥���<�d���)2_������d����Rj��e!�m��������/?,��s��br��z��TAK-?��9�hvC�W&��k�j.�w`I�G��	�ؗ�e��}xWj��(�2Ey~����o��d���N3���u���,�F�J��q�e�dBR��5�5��D� ����J��>�Z��R�ߠ��N����+�H��cܯ�I�=��X`�l	��D�Q�?���q��=VG�y\I�;A����g���W��v,��O8���"[�7����H,�IU�>����U�i���]Ͷk�GZ��VHV:���G�ʄB��DzlBu*�����*��QW�OЃ�tL���|Kߖ%�r7�z��Lau!싀-�(.���o�<�U/xY��*�n�k���ޫ�l�Ю���Zz���T+c� D��0;�+��d���R�	�DT�ϫr���b�Bl��1���%B��h����v���*��~��	�f9�=INTz���V��'��V�˺�i��eGY�2�<i=*Ue���)��TW�c��ֽV��F{�I�ڰoe�����X�`�(U�mHe�d�t�-���.MhD [�8z0�8������>\�'*����p�=Ӽ�[ �+Hnu��F��C�j��^��OܣP��u �U�q��2���a���V5
XW�h_%ȡ�I�daG >Q<�B��~�x��|�_��4U�+U4=���sK�j>u�1�0�J�N��r�W�a]��q�X��E����L��C�#�����P�:���ɰ�\X�`�١�㰈���Ʊ��~Qe.�7�[���@�y�av�;-9a���e䉉�LOp�]��;�A�mC��X
`�A�8������~-1.�Mc)n���:�#�98!�#rʖU��|��%MQ��!R��˒Z�
.��dʬ"�{��j������}5B��23j���/�^{S�.Bi�'���VR�������(n�M�[���V����H@	�Y+!���z����h�"���oӀ�DAv���W���M����%�c��a������k�����8���\��ln3Kz��*�ȐnD�j��M�>�1ͧ�7tl�5��F�d���{	�3L���>��<'<03k�r��Rt�C�/��3�p[���+d�ss�R8)�إ�8�=0,	���,Y�i¡�g1���������}���x���(I�,Ĩ��P��7�s���Η��I�Fdds�m��'�km�����'��Ck���tb������Z!ּ��2݄���(�p|�SI�Ϧ��/е�OΆ�m��R!��Ǌa	�~c*���7��wp�E�吝�;�B��t���XN��f�as䭕"+�Yg�ޡ�e��vgi��S%І����-8!�>>��yYQ��!��e����~&����G��d3@����\A�w���=#�>M�zsS[.����e�}g�pl��P�ZMd��p��B,ӣ�w�Q�X���1���S�^��q�$�H_S��lv1�~A��L<=)p/����\I�U�]�Ԅ�{��Sq�4��|Uİ]k���`� z�M��Z�����A�>��	��kx-X���y�<nse�:��9%S�M�����'�=�y��W����r�_�̪"6	�Y�kp� ����G'�15����ԙ#p�yGK ЋGj�А\�&a��/r�k#!��Ȋ@��7��E��u���~*�� �T�i���ܽ��z�ts���Xz��B��;��=A �Q��,����d�xV]��
���^���#��~�>�(ձ]�g[H%�p�&�އ���� �
����/a��}������)���J��Ύ�!㪽�v4�#��Ƀ@n���v_}�*�z�gXYv"���n���M�z48�Qc��Y��?K�m
bE��#Ne$��k�� =���)qȮ�a��B�Lh����������8�K�e��p.����);�ޣ�_�r�{-_��6d�N���.���Pa�ƽ�'��}�/c	�|���U2��80{�8������|�D�I��RU�`\�&}:EH*j�w��m0~cj��$a���X`��S���\��+�B��$���{�2I�q����S��{�0��I���x��0���>�9;��97���#Ji�q�����{�y���Wb��k�&S#Q��y�2��&�9'~�#��BkO�Wa��!�Y'a�d��oG<�a}$��Z���ͤ<t�R{C��{=�?n=O���ӻ-�C⋚&��h��Õ�q7�9:���̶�퇂`��9+��.;�n'�@FR�pj���Ɉ��]�K�@r�ښ����6��Tx�t� 1��C"K�.+s��oZ���CqC��n/�G�!jl8���/�Y�+o�O�Vi6��Q�Kp�pm�Z?AYm�z�),��	(���M�P1ݨk[L�.ߋR�4��{w�\v����̌���U�g�s�9���J3۾���$�������V�Xd��&�fq�[c�4OdR6;�A�<�/���vҊ=��rr��<nc�`� ��[�	�A���r?�P���rw�.�h{X;W|������s_��y��v�W�A\��d��\�+��&F�S*��r��E]%2�����`��@���8��2%��'kvAyRRs@�d+�Ҍ@ �,~��1x�a7N��G��땿��̣v��Т��v��}��`xL���x�~�.����0�{�.���%�N	�a��o^��te��H7���5|
s_�`-PǬ�;���PRNl8����#S�C�,�_��xquQ�gk�ܜ�x�#:Z+��\����w�m��P��܋��`e��Z��4_��*8�(�$����?��ϰǌ��B?7q3�Y`ߝ�;Ѣ�k��8���Ε��r�e�C%ʼ�0�m��D>�s�vV�k�nD\v��W�}2~�r�{�[.wn�j�5�.�g�x@O��?�|$�t�u�"'l��q�y_!z��y׍��u�]&�<����=| ��ΑQSo���]O�Q��{~u"�x�9So�&���BE��-���'+�e��6H!����_'F�4B��<����:Q1r �GZ�\{�v�����������9!̓R�!]n
X}�@�Fdl�U�W/[gnOԗg_^Tx�a�D�o�I����i1����Ua0��޿��N�R��&��f����ȩ~��q׺�ڼ�/�zϷ��o��o-�ǈ`� <�[�Rgp�r2)�bLmꌉ���8맮}�.�D7�B|	��ى6fI���5��O���������F3��꼱����%Q��i!5��V�5V���"�����q��&�ag{�N-a�#�����%A	�g���
)�ᖺIh"�v�D���l�P�T��{��`����_����gx`=X|v��a�"(k'��G^{j<�r</�a��ܩ�F���:�K2�+@�+P�O�S~��Ǜ��2'�fs�Rm���p��q�� J���&2o2�=�5�}25~�+��U�����M��!��m�D�4��<�ڪ����*��ʘ`��s��܄y�������t�_F �]�9!��$��������^���V����F��n�.�ӿ<��`+ߙm�H:��oA�J����@�z���ː�*��eꯙ:�`*ƆG�Ɯ�)����� d0��� Î��*F�]A#Mo8B�N��� �1\p���-Ʊ�?J�OݨǠ��zbj�)!�/|Qy����n���`6��2�����+���E�A���)�Dl��V9+^�fH�>�]-����-K��:%�Aҵ��d�!*g���;<�C��T��AY��_�����Z���=�����ľ4 ��;#I;��D[xEYz�Έ\b奔�L�s�{�ǖ��?��b�A6�~&|:R �1(���a�34�E������k~�ZG�<�ٮ~D�M����[�a��*�{ �
���
�5��O9�
�|���h�{����2��A0�]��@��F~��Λ��h�S�=�B�ؾLK��7���dJ[��ȕ�s�k{x�Fr��=��}1 ���<�+h�o�r�7����Uq���d���6f�BMל�xI��x�Z�`�j�T��|oq�vWcYvCh�(E�5��Z-DU���m�>���r�b3�#G������,k-���9������[�M�S�Q�r�Q�y�(k#؄hmW���K�~'i���5ܡ�O}���a������X���Cj%�-�p�y�o%��h�'P����Sd��JCу@��2ճڴ+�d�����Q�T�0�?%��.e��7s\�9I�F��RHO�G�q�]~>�z#ha3�^��b�����=����!5�V�D�3�����$h�Ф0V���9!vGś*�;�U��u�-���o�3:;���yO4�B�ȘAȴ���{G(rd}�Ƥ����s5O��^|�[��G*`��ԯ�e33�G���ʕ.��}��q����G����%b/�>R�c���sB�`�A�Ǒ��|�D�(y�bq�=ҽ7d���Y�Mr��Kȴ֏~��~/�q�A���z�B	�"�2�{i�[)/>�Ho�Ќ}$����5V%��&��_�lq"��*�y�w"���I�%�h��g�B8�D���Q�&} ׯ���c �W�rop
}��\�U���zZ��{�0���N�d��%�ըG4j��=5�F־��q؇N�0������ʪ�?��K6f��D���wt����W:O]a�b2��?�ܙ��ߒM��>�|S��;�Zi �C�Ѫ�����g���T'A��+� z��\�5����ݒ�c�}ý�Yo�,�z�]�z^��ي�HZ��G�?'���EәRz�]V��Vc�H���%L��w�Z^�ͥڱ�$��}��n�F�9���k:�Ċ�&Mj��́���0�gǏ�.�0W�pW'���إ��Az��6���Xvpe:v`h�D}]��=r������������{����j��yd�q)�ϽWm|y�.����EF���F0��xӋ��p_?8k$.����"���2�2�0,�*��G-
rB�v��I�n�&<C� ,����[�.a�'�����ӣ+����l߉6������TE7�x*����>�V�SP�D�/�T�D�H6���������R��\��k�X[�_?r�pd"O��a���K6��|���q���E��S�,�����G�=?$e��l��gJ����8ͧ� 2��<����,I��/�Np�,{6�IE^�vSx����,�' ��,��� ���Zb�B��3|��`�ur�+J���t�%S=������Jٲ:e����Շ�|�����u)k�N@��kV֫t_z�e�x����8���h�=�7�M����'5 XV�U*��Z@��f8��"�H�8����V���}��n���͎P�7�mgtX��ޖ���4�}gB�"m��Iݟ�
��2�V,ȩƎ`x�r��lݦ�([�����t�E�����w����R�������`;R3�B��|6%��9��^�7�=ԭ�(���n����R�s�+s���0�Ji� ��M&wRG���)[���۩뻒)�b�A厷Lh��i�`.�~dY��n^�3�o���q�� �$*�2\Nr�xo�Q�hoT�lKE���X��1D��Nj;���G�����TmB��Z�U��ʗ����?[�9'�9��$�:�!`�l�
�.���5p_�l��Y CZoP,v_�=x�����y���v��}��'�ʪ�I����A��S����]�۷��L�Us�np�O�T.�r�Wy���4J���O��
3g�p�*�A6V�1�_�������	�����t����޾��6߆U���B���TN-s�� <��'^]��Pp���|� ����zN��4�^�1d[�}aQ2����~6�µ�m�_9��~�m����Y[<��^\���h�x�'!oj��G��ߞ7b���-b�%贮�-0)�i`��ʳt� �WmT��V�aO��.�̝��(���\�luY��8X�6l����c�w<%~$�����QR>P���fD��Q��-���R���Na�oϝ�����X&��f�D��XGС��M:��e<�Y�Ѵj��h��	���l#�Hc5_�1r]��(�4��k\j�?#�Yr�6bJ4�A�C��)���;?3P��"�cj���R��RO�cL��;]Y]��M�2htӷY�8v8}���(�`�n]S�LyQ��ґdiwo�N�w��#>=7�d7�7Q�p���# ��H���'No��Iw_q��&���i?L���[r�O��-S�muɖK~�7Z�i��f�+}�״����:�j��K~�g�o��c��$t�/ҝ�>�8N���?�1������z��*�Al5%�u7�~��$ƞ���9{]�碣������{�_ly��������}��Sq���0/��nz��"%��<fƗf�7Jf����'I-�o�0E2�KPlVN�CG��\�вo ����tq0�%E�L��J�:Q�i|��5��f��CQ����"	K#���Pě�
d�+xq�C�ϋ���Y,8UZ��:�
v��]H��2�䩺9.*��.#����>M"6�)OU��I\ ��氧��7�D����Bs4?���]ߋ��6ռ!s�ph����-���*Q�����`��@��j��fH�?2��Wm�j��g��#-Q��
>�.s�O����d�Of�5�W��؜d2��
���JD)$�aPV���Y��lo�eOU_�a/F��p���,��]��������y8L�5�&>OK�̎3�!�;Q��@�a�x���GgE"d��TT�	~)�U�2��h[q���H^�ٕ���=�-`��͓B��<�����9[d �3>�Yi��L��Խ�UiG�Ɇ/�$��(q�*~���+�wo��)�_��"Pikw��zC������/��M���SfA�ee�F.0�KpUn�C�)��K�|�{��W��X�u���F�i�
�_X�/9�!Lk��ц&�hz2oh��OĤ�C��{uo6��B��?ƈ�͂��n��b�Hf�Y���QB�X*�͠8�݅c�[kO�8�&Ƙ�>��] q�:!���)ް��9z遊�����/�%��&�:d�VB[oA�
��*.���K�}�$B�9�(<���ʳ��G?�PN繵�>���!��E@� �Sf�ё`���im��K�n?[����Oj)�����h��5��|������#���VrQ�� 	�%�Ht�e_t����8P>�����X{0��u	��X�����bQ��t>��b0�N���t'{^N9���-]5�VA�1貸m	e�����h���t��ϛ^��7�8�C�%t*Y�y�S#"&dA*�Ν�i�����ʺN8��jDv�$Z��t�������п�_�B��֌.��U�:Jg�R{�ۂ���m��d�K�c*�7�g��4Ք�E�B��u���F��C"�����3�کDyj��	�-���.y�w�r��z(�t�!�X��@�� �tr�ʁ"�y��iQr������S��C��������ە�@|��c���bl>ι�Y���)�
���vQJ"�����r+����{����8l�Q��T�m�K�/[�-����7�a>��&���E�YH�M�)�C�`']�PW�-�,�#�������[b�X�:}b�G���c,�0�;�ۃ�Pz�����9s���y@[Im-��dsY��Xb{�΃:ݧ��F�r�EB�o�_u-)sV�k�E���	��E��ŤjI��b�+��P)nf�]s��*RQb�g��	嫎��"�7y6�e2����Uq��YYP%�=&⨿L,e�tޏ��A@�U�6Ja������I2� ]�3 ��L�p��̌z����E\pv6�l�����:��n�� �'���1ّx���׃6�VҸt����0�����<\��`݈�K�R�Pá�2�!���K���mNת4�ǥ7T����Ȧ�#�7��	�s�w������-���\'��O�l�������NU�������@��<c�<��WD�qJq�
�R��.��2������q����H{����b���ߪ��ФH2����%8�͚H"�'R��=v����/�� ��3���n�xC�[��0���uG�8�J\2�ᠣa�\a��މ�1�W�����ӟ>���zz��j$X�.�vOs
�A߄��r��Il���K�1sv���ӹ�0���x*0���Ņ�(�o��=ť6s�m���p�"�����Iq��'��!|�y��B9	���V4��Z�AJ��$��/m�!_�l@���B4ݔ2,����8���8I^���zQ^�l�	(� >��K'�K!�j��Y��j��AE؈��^����"��|K��y&P$Ĩy�`-�b^!(�p�X��{�`s�K��~�з8�"C7���J>s�&RY~F��T�q�����'೦�Ԭxm�ϖ�{i�'�ax�5�� x�"oV�YQ����)/a�f�1�L���N���~�
?oK{)$W[������b+V5�N��s3�Е^H�
�P�:g��m.�&�0:JnA��!!�87ͻ����N����h�>��/��/р���Ϫ2�h��z��wEg$�n��Pk�ݓ:-��ga�!� �����#���'�C��x],���z��%���;7*��$���{$
c��52��iBߙ�Yk�gӱ9��ȯ_�D��*H�sv���5��cD0� ��ÌS�Y�C�yv#c��*��N�d�~|<c���r�Ei��ǉ{�<_'#�l������ܐ-T�@��=3}�Lvɳ�"v��
�кX!�hyeHI9�%���D���=͞�2�ڎ�h}�o�%ϋf��x$�����}�O
�^�I9�mۘ	��p��p+����<�eCNy'ѕ��4DS���*~+�Pb�����4%��۹�P��B=K'��,���c1��i�s[� i�`�4�M�x�kA��Q�zy�4K�f�E3�d�b�wn
fUJYZ�سH�Z҇�����9GK�K�qM�4: PW��������OҸ5�]>#��:�5�u7�xc��A?�$'�&����\Տ"U��ȧ���cl���|���q������*�xjćQ�C��q:n�O7+F�kRx�+���$'�;p�
�)��A���b(oR�,+io�4��<���o���o~��ϙx	z��+�#���C� �-%}-�s�<��һ����R������`5̮���O)I��q>��\�F��2�%JJd��J�!��T~����~�q�^Q�2H�G�]��>�o��SAn�P��k�����9^u�!;w�BZϢ�a��xJ�d`}�|:~^I�m�l�7;��ڨ`��/�f���u�p.9 ��h�[\��]T��< 2jG�RӌNu1=��^��4r,	��wY���k��֞V����cI-�"uuL�(2U5u59>�z�pB��z��@|��fd��*�tHS����R؍s&	��`�����ߚ�>գ>	C���L�������RƂq�>�?˧��4+rE��=�ZÁ�Q���1ۈ�;]qo���|��C�)���&{%��l���|��ж�cH"�)
�l�0�q�u-{�I�������u�y0���7}Q�7���"��>:�L�t��^�u�;��n�}^��@�;��"΍U-�J�$Z�?��4���NT����������4��E�-�����6�k���LTk��x;�s�S�mb����Q�K����/}��J�n8F<�o�\!����t�fm��M̫�5��LD�[G�����*K��=$��q�V3��9Փp@,XK(������ M�.�)��r�`�6W��x'�Z(�w1���`8_��D�d��)�-��F+N��K��R�x��� �7	�0a�O��Ǌ�����P���9s�%�Dl�@��+���̰�@6��.�`�l��.� �!�-	j�A�︿>/?��;��[�t�a�jEv�"�.�ȳF�_c�R�,Z�4Rt��*X~ǁ8��?�ٲ�'b�gN1��R�t�c���ӢXw��c�C�3ƝڧkA����6v q|V�
 ���*��U����V�
��g��9r�W�IG��5�a!��U9}�g�j��ǻ�,P�zK�2�����b�V��tRN�t�4�PG�y���s%3v5�QP*5�'��;�e��I*l��:+!/�˗�J4�f^:e��d��ͧ �x����fB?5��C�
u��n4JRg݋M���.��Y
6͒����u�.LH�C^�r��+���
d�mB�g`�>��H�C'�����9��:� |� -��,*�B��O_U���b�F�����ud%����f
�iH�1uS�0C����#��_�k��Z,�Ϥ�|��]�xo�h�i�~����ډ�W,���?��I�%H_|��׍�i�=k���ӳc��d��7]@��v�E9?�1PjWE�lێ`�Xx�?:v���s*Q���Z31����WkT���F��T�f�S��g�]��;��p1fc���4'�#����6�ix��S�p�%8�@��e��7?# �K�e�4J���w3��\���Сy�1L�TmVW0��jJ��HsЉ �8�`�xu��7�|�%����G?��@a?��劗iG?j���x ���Nə���	�Et'�s��y
A�dדŰ)�4� F�#�}�<��c�W$������'��R�~��Ċ;���BO�U�Q�F����5�y�Ħc:_7�/q�|Uv~���:M��<d�䵭��� �R�|=Mg�͇�>�·a�b�'�	��4���'&Y�j���ʌ/+ǔN��ϊ��	�u�]V����zG��V%")ՂqJ�+A�#�	�Bc7ɔwqҤ�E!&6�E��õ�h�֒z@Mgj�W���:���n5��@I��jm�E���i�ϧS6E[�K�ҙ����j0��!�2��3�e㱺��z<�D,��aȣLWÜ\���6rަ���fF9R<��-7��oQ-W�c�6`��>ܛ�8�$�~iX�
wba
�K�N���ߡ�����پI�q��}��pb9_�����AI����aUD�t(s�k_�ww��Fۀ�>�V5���	�2�J���+K��Θ��6_�"�ݯ��*O�*;�T�v�T�io��=���v	����0ƜXav�_��[��+_5P�������"���`�n�����=$H8�
e˔(�� �;�������O_U�d�e�D��2�M�b*�y��p;8
����k�Av�ϲ�����"���z]��W�u�U���n �g]e9����=�MN��r���s����>z�>i}F.ZtV귵�$pb:֖�CРaI�@i��d�A�k�l���������Q�bF�jO�Kɦ�S��:LX%�@C���_ɰc!s�yw�!�f���F�_�-�#�G� mؓ%��#Bj´��<�q�L�)��¤YFȭ� _��-�᷈�y�H	�ˠo��� qIv ��{����I"+V���2~��M��q+�A?~���@1�9Y�j��v����N�(ȠߘZ�ڗ��!����z��.����r!I���V��9NF��)F�A�1��c[�:�Q�)�c7z�S��2��,M��-9�cY ��d�ܣ�-��h}}?&F���V	hp�f��3�!������:�U�p�Ҁ���'��2Q��B���Ђ<	�gq��rw���*d<�I��y���������~G~�Gʷ}�J��Qx|�t��ŵ*d���g���8�'w���>K�{�u���K�i�|���I5�4�S�ڸ��w��VY/A��x/u[9��e�
1���YD���ǿ�-f|9��沈"��G
YmLĹ�9���)��ݻ䞻��)�
ש?gINyh�&q6�D�t�	l#�X�v�:������)޸\�g\�|�0�Xo���:\��S���dY7���{����U*� Y��tZ�TҌG�r6�䞔)(+�%�����΂H��|'*m�p�k��.LQ���֓�y�Q{ķ�'yqfc��������y��O	��������u����ҕ���2(�'k| �m����'�b�(�&�%Q��8_�T�����N:�u��05RTl�8��A��G+�������~��>����W�FQ=0��7�7��wj��+�`n�����.'ґ��ޣ�̈\C��!���](�5��Ed�I�'շ��moyp����s���8P�]�`��J�j�`�u0���W�7�{�p����	Q�{.��� �I)��Ɵ78q�/|٫���r\��qu%Kv��3r}�d���_^����m�9/Ⴐ4�\K��\���+�c&s��`E*�6��+=�P(�³��ǟ�1�i?A����StmS��OD�����̎o����כ�}'�+�Q�������1dR\�`F��g3Ӆ1�O摬�g����?�ra�h���I�ܚc��xu=Գ�f[\��D#p�� ��������MwFB���M��*m��H�A��%�l�.�GGf��qx\q�0"��&��E���"r�i1	@�Gÿ�
��֊�Z��7��hp�Jq�"a�1�X%nc�[n:ȏQp�~u�Y�s�'z�d�U�$�i��p��NK�W�/��n��E6�����7U��]�R�ͽ��I����û2��)���`���.�l(�<���R`��a�Fq	j]?���n/xp���rVĵ�µK���O����m�+��>`��c{�#E�$��xH�~)�m���z��y���?c�4ͥ&l�p�+8��SG@��u����Ish���st-�?�	�g�GGR�O�А���q�-�c�5kyIV@�O�;�)�p�Nf/��7u����A%�B���>�be�5w�J�Ϡ��v mA���Er��"�5qW'�ɲD~���X����&O/j^4-��*�5�����PX{��9',�:-U�nK��V�v���
v"��2+x��r�Zc���åT�ҟ��&Ko�:Ag�jT����2�^�`�2�Zb���{*�������@?���$(`�ݸr�2zt�XbD_Yqk�FE�f�15��셌x	�-�֍}�m	5�dR���FPմ��D�du3�W�Yb(݌.]��kI�z�(���TBKa��������4�Toz��t+ i��qJ�AΫ �����<ٖu�b]~h��o��4�ۊ\Qp���d6��ڙ:T?�C?�j�y�H���Cz�=e��|pE����g���7Bp��.�9_f�b��1��HC�����,Wn	��X�/Oݫ��e�0vm�s'����.~�3MMc��H�2'���c fd�w���qcC�l6b�gB[N1��x�t�>I�Md�2j�گ���*�H�[��p�Ti3ddRi~��ӌ�VL֤��)�>ϑK�?0��\)%�#�a��LJ���0��[���ݠ�uo�J�;���1�D]�����	gJ��c�^�3��Smo)�m¾ҚQEh�z�z6P�v�C�v����>�'��EGF8��3��
��G�E���}�����%K�z�b��Ȱ�B�4zs�,��DV����S����E��Wm��M/'��h2����yʄ�C�c$w��KR�n�_�_�u���!�꺪�)�x4^kFۘ4����`�2��P����e9L�zm��P�s�|<��s���{cO �?;���;��7Iƹa7�sh>��t~a���M�������<��g��E�#�vi@�Y���c�)5�t��P�{��r���1}�v�B���O��Ws+�Y��ܫ�3Qv[�õ����݄��� >�m�@�m?�A�l��z���є�^v�E�����X�pl�P�>����ksI87wL�75hh�1���ؕj���0aR�4/o�7��0C��|���3z^�+�~�<bۋ�D��)�~��A.���{�GH̺Yd�mZ+��G��.m�2��]�!ǊorMU���C�&�zU{����Th��oH/���$3��vY��W��S��O��m�>���F2���~*�3�>��+���c��!J�:�>�7k��4�UI�1�X��n���N��$�b�tJ�Es7��C�C�n[^�O�2b&|��mt�[e�1�f���hEA8�6x�X�q��*�m<jЪ�^6wj0��S���2�<=��!`>�$m��6y�������3���2{s�4��%��t`I�z�lQl #���n��:0�)i�@U�}�"r����Ux)x��b>��i��,��=yaȢ�
��yJ���&X���v�VG�О�G)x�?@,�>�'$ˊ��/��I3�a����͟E�;vc��A ����͚T};��ң�L�:7-~�6Jm�g���o^!�zX_Rv�L����u4����4�o�����r{
��5>���4�����P�=Ҏ��[���Nw0a����r�{2�a�rz�-L�	��1�YB�O{)����ޅSa�m�x��W���b��%�;렫}=6���m(���*�����5F�n��S��e����vINv���{�_*so�J�o�m�o}�8�rn�2��l���\i��à-�������8T�!O0ʇ��	��(m{;�������� ҂n?����V�(�0�e�����~E�� Y�6d��E����a"�{P�J�m4#j6B�v|A͈_a=!2�M݉�U��<.�)����<p�a�0����6O��KM�Vǵ����u�ˡ���,������ٔ�2��l𔳻q��fϐ�����ږN+��"��Y'u��B��+�4��6I,�Xۂt2�f�0�7�p�[��7��w~v����₊�n"�4��>d��u �q c��HqT\�׹�0��rkլ���#VP�]< ��]�B�TsS�&�F�SN����:|�h�r���m��o/����n���c�#�0k�K��;�&����4y%�2�L�K�Yw��p�r�wY��(�:�l<�A����xM������̉�p�d Л,���k����I�t��A��s�f|��y���|I��L���u����� tk�cC+�Ɵ��~O��,�+�*s�&��粁��L�!RS�.�/���ý+�Um��([zי'ɰnu������?���-�g~8&JԠ�ă�%��YH$+�(%u����V�C���в�	��QbQ�۳5���7[F���+��	%+��0ܬV%�mӃ��Emm|�1���#�iOz7yU���y'ʓ��ϏM;�.���[`ySJE��<>��İ�S�K�Q��e��*St��1�Em^�D�X~�d1=N�!�2�e��:��y����IK#ӏ�a���֝��,ѵ�{ړ���|�j�N�� -�)���l�v'��|b�Xx�l��497�����;
;2����������k�ȧ~D{��7��$WW�p�j6yѐ���B!��j���}�@~5^�Z_ڗߧ��t,ǢF�ɪ�	���ly{8���]�E@�U�^6 ��K%q�\�AH1n�����hm�\~'"0?�a�3ү%��d�����P�m�HϿ���T!/�ը��F�;�Kta��Z�}��՜�pih�%��#��wy��NX$���e�B�c'�����zCU�Ԣcb[Rt����v�+oF�y����R��L܍�|#�
��,ez
�������٪ćH pL����1�^}���ˀ��H5�^�s�S(*eq��r�1M I��As8�(�-�<�q��@�/X���A/z���''d\�J
t@��]�`9�}��7u��73�D�r�c��-= %z����"CfF����SO��`���w����ɱ�X¼=�m����_{`�L`) ��7bU�NL{�s|��I�7�-�-�}}���9�4� �v��]��jX��t�v�J�v_ї.lΔͰ`��)(<���Z��i���sP�Ʉ���#�$��� ����k!�&Qu3���:vh��詛�_�����w�cS��Rʊ�e�-��(�w�Y6lu�R6��땩����Z�m?��h>Z��yq�Ynj!��\�����Ѝ���V읁��|���ghC�I���Y�j�^Z�H<b����o�xͭ�K��B24Y����u������7ypgA�У��dM��k�s�X���f��=�d�)9��V[gR��!W17OTB�ų͢č*�B��8�CK�)y�`�~|Wv�1B"��7�J��͞����f�-�.GG�a&�3��-�%]i�t)�,�-)�0r�<�cw�h�T�Y��9�Ѯ)�3����n�{�,ܾ�6a���f�f( zASB6I���|��1Gu飘VO����-�^\R���lv|f��)�����j(��ϐ����Bho��-.����qӑM�K'�(@�*��u�WP!�[�Q=9���ڹ���)N%�i�~xzWB��H���C.�43�_�wȁ?�,2�|Y-���dIF�lx�����#%��'2���k�1D�����Ԇl/��m�rkz��&�-i>kߋ�
Hry��Ư����;�|�����s�>7ۛS����{*�*b��)Zh��U�f����o��g�ߛ*�����p������*���3lD�?)��~�#fT0{rW��Wj�4-��/v�v&��_z"�/.�cn}��!4H�N��3-� p"���LmU�`#����b*����\��
���r'���^/{��b����˱"w]�}��2����or y�>�w����n�_��UA��v<��hڤ�x��a+R�3N��pp_�7�hz��ŵ6�''���2�"�M,���w��P�bl�3��#�%b�;���.8�Zu���!��i�"�<˦��C�X�G���*�8�)��i���[�Ě:�{[
�?�y�*N#�z���^�D�aX[{%�h������HsE]o1���9 �F�߻��`MZ�`��Q����+wÞ:w������B,pa@G_����X�sm^�6�(���n�g��f鳎ɸ�X���(Cڝgo��V]�2�)����=�[$E�������X՘"�˟F	T���B�o`^�QD'w��aέ9�-C�E�x�-!���
���,"�	u��C��қ��8(�K�M�w�z��$5[.1s�ʻ֒.�ԋ&�����߅�s�˪u�<�����l��t!�ԭ1Íf�x�,�ہz8T�d�D{���f�V��G�L��Dc�e�|%h���͚F�_�\���:�b����;�!a���Q����z�k�F�Y�r����c)�Z���Р"�'|�s���E/����{CҌ��N,��=����n�g*����<+SQ��rP��H�΋:l]�=�B�|�Q�\`�J�Ջ��=<��ĸ�l��<�z�Ê�VIe�_��L�M�{y�H�b�$t���і�x->�Q�o�a�!nѨlS��Ռ��^Y�V�)ݠ�>�E�ڞ�ڴ�	=�t��Ғv���o� �e-�$5���;,|c������CW�ľ�����3�K����=ŗG-��FUy�*Je��RJ�Q�����|z���ҎXΤ��Em)�V�PWS�n�iɪS�y.U�ŷ�5ˌkQی���=ji��*�uTy�J|&�`�p�+v�7�����pF����;�l�H��v�y���;GN�����$NϞ~G�U�!5��35���h&���9�9��X�1��`ǒ��IΕo�َ�Z3���	@cH �0�!�*�#VӰ�m_�]/��:OM�JH�5���ŴE��Ct�w�[6��H(>�1�@@�,�B�X)?K���	�ofR��d�t��#�dF�7z�?G=��y��P�u�~�ҸΙ��@_`�=�I��bq���g6��d��AnK���;����E�r�n�w�z�/uT,�L1}f:*/T�}����C�DQT���nD�"{�haQ�Q4�^�i��#yl}�	g�֜�2��x\���"���A0�%��u���ue8v[�+�4�ZC��&��x���ʷ1�_~˳�bH����~ڐ�?�?���X���q�y����I<�oT$����3@Y���1��O�$qTs55fOf�˘Z�&�CȋhS��yEi�:]�\�O�}�:���=F!eu��o'�*l��Ѯx~��NNW��k�]f_�a���ڹ�D�^�G鰺��T<��࣢,��x�%)>���f	7�K��Y�hL�˻�E��׳+`$apuf4b��;�&~�@3J̽f�D�fm�pl�)� 2�⢧��U�Mv&.��ؗ���)$�:����R
0  ���E%���$��k���"m��x2�������S��""��g^�@Ф�b
��)[F���7M#9T`qޛ���R/�&r�\�O
P�c��e��O����f(p0��nS8��V����WN}��C`?�g��,�=���B�;�M��k�v���
�y�;8�j�y�ݹ~�)ds��RSЦ�^Ъ�[%Wbkf:A#$%���^���mkP/�P3{1󆮲��Ok�	T�3:�@r�yX�Ҏ�E�V�@A ]
>�R+7:�0mj=h����'6���b$�'`T�m=<Z�'�v&@p�i2Oq�8�����4��V`#[�m
�����kvjl�~U��5ё��kP�	`"��,��IrW��d����2��6��eW��$�%���FgVh�LBb��H�h�e";�E�OT�@KZD�8hF���Yl���ˡ[�
��g�˟5����7j߿��D)�3��Ft`�-�5���>bB�C�M�E��(99UU�J-ޗ.�%}YHb�>꼰&M�a��m�Jhp�c�Y�ߔ�/UO�P�S4iؚ�MlL�%���=Q7���p��o�y7����Ln_�����6z7F��t�;��(�֮��v !=�`?�j-�9.t'�|G��ʞ�ǭ�{W�o@<L��l����$�K����C�(��	��Hr�뾠/��� � j����l�Ϧ�=3�m_��ׂ�f������N����F�w7ӗ��n�q(����gI��v3.���;�<F��|NH�T�.���.����"]�����[�S4L���D�Y�[p�3��0�X����h��UJ3.*�l�j3&z�r�V���þ�%�'�}�����LD�ؿsŁ,�/��>NUE '�~}�M��u���H��������������$!��&�3��m 7�dt���� ;CY4�/�'�+��_�c�mcrz����zxYxC�:����ڳc��ncnBqHC�8�Ʉ�f/�q����*��	(+7hbͣ���e��A}��vp#��Cf3�<XB��=J���>���� $h��9V
ϋ�_��9�u#�C;9�d$�<�����"V�Q�b���k�
�XSgݯD���+R:��e݉�jܾ�Κ�X�O�̰hmI_{��|��
����aXxPP�UϦmlӑs�%�/��%����g��7�$�����)�6T��R[X����T� �q���<~U���:`F��;y���Bv&���xł�iI%���R���O-*�IV�e�B���p�稬�ݓ)�ŗI"��i�\D#�t�{.XB ��-��X��2|&���J$����$�1+<��㿯�d�V5�lt�-�iǘ��s̿��)�$��R�^_TN3t��U	<��rϳ�4�r�^��u�T��Y�ZՈ@��i �-U;�#�aZD�i��Z_b_<m)�'��5�,��dO���\�0]�i���{ܡ4Y~�W� *����Q:�o�W_R�4���I��"G����,��
X҅���6�j�sY�(:6��a���=��'���=�����̨5��H·:�j�@���W�g��Hߋ��c�Z:�ڀ�o�\���!�;�m>��3�ş�0yH��xfّ`�vnN�i��rjM�)���Sm���򫶬��:��є�4�@���&�i{��Ij5�˳�	�s��>��x/�B�/�{��y���F\���X��t  _��9�ꑦ7��K�Ó�ƪW�<=�&n	�9�����ZAV�%��1��Pf���SE���Sݝ�����w���������XVq�eRC�h$�AA��t��t7J�8�M��h�����z�G�'AF�����mD!dv6Η5�1�"��K|�mdeR�bM�5oFn6G�+���+'�Z&�Jnℝ�}ZD���	M�-OI��Z��~���inCp�I	 �Ş0����~fuJ7���ĥ�<m�/}�"U��dQAfUYJ�չMP���  M\�u�������(.d>|uFۿ3�ζ�}��w�Ǌ�P�0�8K��[�A�ɑ����J ��Љ��,�f��l���"�F9Ox.�ˀ�j�d�h	��%膎e�/��#���ʛ��P���)�z$B8������2]�n����\,>�I���C����r�#��+ �[H8pkxy�wH���m�(��B'w�����J��#�>;�/Y�;-e�V���Mڕ����q~����w��Á!�G:!}��5��sU�8��`ga?Ȇ��Җ`u��&Q� ��
^I��{o�6p�Dt��_��|��>��~�]���4�.�}S)Ḅ�A�	������n�\Fe)kuo�V�5=g6��� ��%����O�ԁ@��5n�V˛���ql��M����*z+w���F��'ՓZĐ�x�ɷw�*[v�=�Lp>ɣ�o�X���A��l�H/"Ġ�LKvR	����.)��X�z'���Ǘ�c�P������hb��j�U8�U��ű&�M��1��ǧ8:>�,T[�P D[�gZ։j���w�ޞm��er�m���c��p��p���vQz����s; D�5g]�gq��)��F�H����>��(�ީ-{Nl�?\d�N`�=���sc	�?�Tn��pk0� TUAE�-�*g��?�6֗PE�f��Eb�x��2^7/vl�,����sHq*�*� �zq�
�zAE�_�茳� ,s�j�܋��}["�J���9�Su+FX^�ˆ-�#�zf�x ��U��.��*��PS6N�s��2�]���I�|�*��=��Y��zF�7E[GMȫ�D���Z��������ſ��ђc7�ޫ��H�7��Qxv��%�RA�Q���ۙ���1��̤Do~"x>�E���9��+q5*W�/H*��
�]�uбazֆQ5f�|�Y�#ߺ�k��W�#r�����A�#�jg'Q�� �C �s�,��s�vZW�`��3�;�����I�YC]bV��a��k��0[<�X��8���^׺Nzy1jZ�9��]�PI�~���gؐ�;gs��E��G~������������"���Q� ��={G��$�s�v� ��.��v���%��C�����P�}��F�F��x��P�*�ý�c�M5m1	őLP�(�*���O�d���$\DQ�w�Ԑ��� ��f����c< �����z��}w���lt�s
�^ťqM�As��f,���gw�l /Lq����IH��K8;3�2����/,��P���rh �&���5U���h{�X��E�$�S�ރ|	�������k�rHâ�|-�B�=C�p)�ܾ�Y�k�Y��o�l&�̧~M<w�/�QkY�(�g~n�(��c�iq+�	�@�U���mW�MǷ
{��ѯ����wW��ߠ7=Nߐ2aIc#�F����;f���B ���e��l�/��Z4��� ���SGEas�V̾�L��]L� #5���'�P���g�z���0H��#���押9��h8˺Wa,x�X��.��=��Nx�Mą�D�X-�/�. k�P���I�D��=�m(L._��銅�	�pO{a6-H}y��lr[~ʴ"�y!3Q@Ժ|��L&�9��L��|C�m��`��u�۽(��ߘ"�<���ew0g?+W�f)�6����1nj�q�j�Z;��C�����>���Y{�Ɂ�r �o$6>�����пyl$Eqj�
���@�_­t��DPq��9�#m�(��jiv>`���-YҞP\�]4�us3$h���Fre*�]NY�7��-Bk��+&[z���[.���
��>��FMĊ?D��˨�w����N�|�k,Ȏ����	��x�I��1���^����^���1s�Z�.Z�(����!�'i\'ݬ�ac���Tq��Dgz,sټԁ�	�3�����CE�J�m���������i���k�+�I�h�\�t���������G��tCN�(��<���1��g�ð�h�BH٪�q����;�g���2�������6�jBG?�%
��6��/%���d+�QY���'z�qx�`M;���k�f�C��$��_��_b}�G�1���0���[�ĥ!��.u�ݴF��M@��*9TЧ��FJ�m��hy����0�s/��X��^S�!0EL{x�tR�j$�����̳߱y���������R��G5�	rp-[�}�[�Վ����/1��?؂��W)���,������-��W?�������^�|U�P@Q/\#�ˬ��.B�%6��Fz�:\}t�����<�IM�H�ߜF���T��p6]���y��}ksD��l��o��Fqn��G�����1��f(���a�%�7b/�Ӊ�Y��t��3Sbc�y��y.��P���OY�q<�4�Ow��bƏ�*��T����o�j�����NI���f�~^�&P����KtvW�P��uBTﹴR����K�[,^�]'<}�6n��`�_���n2i:���1�Ҕ�t΂����,j��b�^0G^��D��8Fr��6�_nٍ׾��r�+�X��N���-���W�æF�4�҉G"w�,@pE��u�ea��԰m��r���A>+'>∡Z)Y��C $"��KWo�3R ���m!��x=��L��1DP���(k(�7o�j�G�&�>6	gVFC�q2�c�:j�o�+~!����(���D���j��ArE�;/�i��x��*�b�w�䮈6d��,_���!9���#}���]2��������pH�9�03�8:�p(� =1D���)��e�u0W9E[-E��Q�L�|��7
Q�LڠTIhS����GjX�J�)΁Y��u�`�d�DA��	v�#5B��Ή_@��c�4�`M�C</��|߮�D�h� V?��;����)�2�+<�	JP��"�Hɳ�y�k=�=Q��a��$�˻W�4���^ς�8��H�`�5*]:<J,�y��8F�({��Zs�9F�w3�v����>��a炇�����q�m�ۜ�5��.�D/$Vv�p�%)3t;Aޓ6w���7J�z"�Qw�HB��~�#%Pdm˨����)�J��8��DlJ2�e�\h����k�(�oq�����>x�ʙ
�m�kc����z�f�=#���to�'�I߸u�qW����>�"(�9�ͻ1j/�0�LwzO��"��g��MTE�ߡ���e�8ٟL��m~�B٤��J�j ���J+���
a���Y����j��p.�y��i�u�sn�'Ie3k��7 ۀ�X���>+�$nr_��
�_K>5d�E40��{�[�݁l��8��b�����K(S���l���?��?��G+�g��I���ݶ���������p���1|�-�~�Sɼ�V����w�',��j�NVn��<�4KsA����nDtWѾ 5#�+�O��S&��R�K����季 ��7ʮ�Pa>��o�L�KUL��,T�����WT)�������lܮ�¤�w࿶s�� �=z�|/��Ă��g�Yk#���;!ڋl�jn�C�bRi�G�I���"��T�	�f���#2���3
���H��}�������V�G<�����|e�2�H��@ބϕ��N]>%�3m\6KOc��=ʤ��S=(v�v�(p�q\m�lh����+j�i��V'���S���G2��1�	%�g�a�O��m>q��X��`�ү�B�N��ݏf2�9�w�[f�C����tf$'�q����)կ����z������i�a�<m$��Mxnϲj;a���s��Y=&=ƫ�9���MZ8��Q;&���:�8pOn����fwҶYXW�K�so������)+�&�c�G�3�TOB�l@R�K�1���jT�P���t0D�DF�v����~��T#.��_v�V �����kr��t�XJ��V��Kh�Z�dB�y��"}K�v����y��r�2}`�3ܸ���誦�c�X|��u�0蜵(z�x_́�q��r��Ѩ�>�RV���Y��E�q��~M���B,Sw��ok�g�����Р�L쑆�ƒ��C"}��;�,�w <؏���<���A����{���Bc���(H�wmy��"�#���o6���ʘf7��Ğ	�Lnh�Q�E:�xD��.��WԸ���b�����dl�Ǌ$��xP�4C�V���T>�+i�C���b�u@���{��9t=>�Ð�h?�Ѭ��=�TL.���<���ǆ�F���s<�1]�}{�T�_��a��
l���F��4���DM%>fJ�t��W @���z0��T�����=./&��V�r��0n�mg4IX�eY��逑���>����ZZ�EI����V~��s�U��
�s��`��aㄸ��a[i�"�'E	U�K0ưKob9T��.�ls�SV��B2z�m'����B�+(<,����+ڟ^��J	��7y�R�J]W���r��܉cjq�A���~�)�G���\z`�m�tس���9�L���4��)�G��
�S�Y݊��:�z�X�+	 �2P��	o��#@�@�rL�����G{?r��|V������ѳ���C`_i?TO�.RX�e��]p�
���u|!�.U��}�&yb��Vg�ܑw����ځ��hn��i�]���Y���|����%���5+�L�%���6�ˍC��2�FD���hW���*�ެ���E�Z���vW��W�9�L������W�l�5!����.7ך����h�1�~�.����M[gg1(]���霺���o �|<�3;@#��%^6�>/���m�U���8|��怕�	���K�\h�
"�A��J3vO������T-X�pt������=�Unjj�ɆKÁ+P<�H�'�\������e47�N�CzJ�<���/G����vʁ����c}�Y��Bg.2��(vqt5xV~�'�R�ͨ�L�W����p􎐶7����m��lm8@�VEp�ͯ�F�u��j�(zл�K0*� �8��.�𲺰|��R�S�@:��[�q̭�'h���C��Հ�)),���LN��0�O`^��2���v�t�v� O̵W�����>
��,����0����1@��<��9�Vku�Z�s��&���:9Ï�c�֠֬K���HJ�?nW��s�$���uEy	}V�V�e t�8�ڂuy�5�^��oBV!�՛G|"�3�}��*��AY��%ʚ�>s�6�Tj>���7�Pu�6o@C��0���*�r�S)�CRw���e�8�n�V�6��Mm�|	�/�ǻ�����Z�mg��CB4�zU����s�I�7Z$ԍ�G�	ZF��i�&�<zT���֝��a0�t�t���{/۫-VG��*��B3�f��jySD{�k�7��Ql�8��b�DͿ�W+�� |w��h+]�Ħ�읏x#���:uX�э<l$�n\�Lr��IEW��G�����2:P�����:�i����d�7�+D-�b��O�J����9VXd�4�O��"��a��B�cR�f� ���M���9Qol�����9Ln����)�X{ɽ���a�
=��գ�B�Vt�`��J���a&� kw�4
suE���P������w�mW�(�ۿ�#�g%_�{�O�T�X�<�sOcJx�x[2E���T:�����tql��g���c�Rˈm�qo�E a�u�񬟡�K��~�g��mQ��<e���~J�r����D�D��Q���QU'qDE�Q�8���vDn]ؖ~8���+�=��)���1V�o1B�Vʓ�7�35ʼ�&}�������M�����M��#��>̰9;O����E$|S5C��Z����@m���&}I�
�@B�N�1Q��#q��c�6C�Y��V	宗[^W4`����:%* �4{@�u8�5ZB�?�;!U�[�7�4����k�Կ�� ��m)k��y��-���N�ާ���b��T�c�CXJC*ʏ�a�}�5���5L�c|si���8�ϘM $6{@����ٺ^��)����C�/+���I� q�����n��_;/ɱ�2��}o?�)���R��D�qTy�Eo"��Hێ�r>��[�2w�cU�JZ������r���^�
���$���td!���HBr4JzG��YĿc�ԅ}�`��V΍�P������W�zo�����>�?���Vl (;����9�C�ǰ��G��D�*��@[��*�A��L��g�>��Pq>:�]ߚg��|W�~��DB���cu �Mͅ������� �#�����GZ��2~|��:'6�d����N���A>6��k�h�L�T�Bͧ蕅�X������4��C!L*_9qE������z*�IRb��{LsO�knn(���Ȟ�DP��P�(���GI�nMNN(s�u�;}X�pA`���'z�ڠ�3��f��o&������\/�f`0���\)���:I�UH�!�����K��o���ǪYx��CQO�UzE��ひ�L�$g���}�i�52�d0m��U`���_*,y`��X����L�0G�	�oTT�N��*��4&��7!S����ǅ{�?���6�cam~d8%L�M8-��-9���[O�Qu/���}��~{�r��p��} �;�m�'#gY�e��()�=We����d�ap*���BE ���P~�b���5��=��ϿP��v0F(�������iTC��ǂ쭱
J9��@<"�=51�����8�T+�=�N��^����}�9��=�.����6Д�7�+gh�tqD�����yR���iO�ҁ�Q��O���Е`��<T����_L��SKz䖥�$�؂Ҍ��aX�R��5�&q�`������>l~�	Z��&C���d��YZ���fg�H�Y5JF��0w�=�7�$�f���TB������5��y����m�q��͈o�#��
�C�Xm�൦3� �b��^�����A���K�7Õ��8�3�t�g33�X��`2�cC���V_�C��寢f�h���I��U���X�-Z"�S�E(�8q����+�Ž�����y����%�-Y(�,���k�'骅��o�z]��b���"Y�m��������ͣI�i>2�>\UHO�~�	g$�Țf{���x�%A.4�������{<?Kħ`{�=����H���@C��S�&���̗����z�%'�b���׼	�sO7nP+l6Ca�J��͏<\�)a�/�i���<��JCB�󆫱�93X�\��-`��
HL-h�}�3C���XP�j��Ӫ��-�~�x�k���'k�!M:��5ȏ��B��嚞U��p��s��9����:�f}Ao�f�k>M�S^�.��&?Py<6�$x]
<��t��=�{��6������[Z�����ẵ�UC@N*������&0���޺���`��QU�s��&_� ̛���7�_�ư÷��WGo�jT,�^!�V��o~p7K�	�Y]{:�w/\��a?�^��1�> ��j�}NJ�ޑGb��IƢ��by�ߊ|��y�@����+��+As�?�5�O67�Q�E%m�Q�����"�����P����sk�d>��!4�
����nl���-��i��N��5)��A�>S&Tvz�1CN# �2��/��#p��.�hP �HlM8ev2�>x] ��=���.�������E����^�%����W��Y��e=�xW��I�/1'Z���A[�����r��7���\��y��j��a@�cI�?�a��֡�`B� ��F���������q9��C�I�\��7�� �a���=m�C�?���!Bs��9���ƞ`͜-޿�We��6?��Z�@�m�W$@�}��'\�6	ֱ���`���&4l��kH�D��Y=�̅�ت�}dנ��>���� 'i
����T|iE"��U����Ր%1S�mڡ�0����0�Hyǃ׼�R�j�>�
F.8���'��k<����-�2�o����8�J�o����a�ˑ0ӗt�a�~���|H"_��Lֶ��q���K���`M�7��Q�V��!�T����}QE	����#A%E��a���eEvߢ�����1��!��q�o��J0ƒ�㬹6T<�ژL'ť���LA����<����%n�H%ZQ�Ǒ��k��f��&EC�C,���!��>q�} �0ǉ�����z(��S�{+^ۋS��)���M��TXI��~�i�y��T��p-nK{Ɠ$�=b�S��WY֜H� �������"]IҩK,V��u��h=�f�iX�^A�A�,��R}���I,Y�^�i���!�{���&*,<<m^ŬJ;�0��0��<��3~�
���n�Ń��H�}teH�����z���̳�E�iz�[���o�i�P�l8&��{\'���k�j��-k�R(Hǋ�s}H��k�������D���")���o9�q+��ϙ��j�����`����%��d>O�x�B��Qi4��d�.�6.�{���A��ւ_�3�.�
"4�<ܙ������*6���H��Tl���v�j{|�PqK^�6�qG�"X^�QF��ϓ�J�`�3b��|�i�T'�+F�ЪSU�׭����~�)��g9U�:G�]��ӫWP��&��A��	�I���uz,L<��������P�v �v儽���k��}j�@}��ŉ�V�y�6��R��B;��M�$�ԈMCܥ03�x��G�r�R���i�S�|c<UȏB���J)@�J������a���vCX�識�Ӻ]���r�rO˿b�>��,D�,�m:�k��cj��~+|J9;��
K��{��З��j�-�_��S6��f�o�yŋ�`�@���$��p���Kҵ=�g�����̅��j6f3����s9#y�o�s/����Ҵ�O�������%Y��ǃH�4p�����*s���3��~�tub6`��o �/|�z�� %�\#*�/{
��%
9�K�T�w�M[X�v���{��ʏ�k/�v���oa��o?O���csʲ݌&�}Z��.��;�ܼ:�~F�'�n
5�(��*7��=c_�uP;<mM����?m� �2x�<ǥ$" ^��"=z)=��YaO�_�-O�:q�6.+E�d(a�m��Y���-]��6	I{
=l���~ ��[��ܘ~T\R����W���Q���C����2�I �<���!A�����y`�ד�u]�DV�K�*�����q�0踕�g�m�6��!
�k)h�.�z̑��&P������$�]:��?��ZM �3���lX������n�����_��0����g��5&�dx$�l|�%i��� �^ߩ�9Ck����3��Uy(w��ܥ: ����� z5=�!��/�ϸ�������[����+`e�1Qy����k61t���MӣW���uz����|�q��p�k1����\�̳?�n�U|-&�1�f�����?< A���摪��{r>�83�H��X�ܫ �w�	}�I[��;��u�/�� \Sz��11 ����45����� ��6��)���d�����)�sd�Vå{)H�S�nT|_���}��U����28�}��������}�)X#laP:	��-��(I����"��4��4�ߐ��)����܎R9et�^��s��MJ)D��JT�8�Xv@r12�@��Ϳ'�鱚"TƄ��C�7W	H!r�2@�����9�ñ���U����S���&�3�"	��\��ّ�[*���>�����9�ӽ8��Wᄽ�6�wn��K\�Ӵf�@��lr�ݛ'�_��Y�50�;��F�B��	S��� ������ �L�/���c���M���/h���'�tZԍ��Y��>�Uf��}
�����fq��'���C�B}�C H?[`��]9Έ����巵FU�1����|IԳ#�1UTWҍ�	�i��D_���*2w"��2������v����)�Cd!	]�w��۫F>f4fn���q�֛ i{An�*�ҳ�6��EC��J��U�q��$�$���SkO��BL	Ǫj��i#���5��gρo��]�o���S����C��{
J�3���B%^��)��X��A�p��CdV�Y��n<����+�U-غ�m�K��n��{��`������n@������8��29�Jv��jV՗Te���<��e
�\c�K�-�	��j-]�3�8AL�����5*Z{���'/o�?nMз��	_�+�a�ҍ��`%��Nh��Ǜ�g�xT���!�������V,r���֒��O����>Ė�����(�e
�0���s��]�'��!�;�e��(�0-QwD��	/�X���Ph�����^MZ&0'+�AN��ޛi	V
?�/��];������nq�Ǧ�|��.Ӎ�lCz�t	$�b�a)va�~�Jq`^$�8�.>溞��E�Ea���
*�G��u�~&�eO3|zҢH�2��(�~��Q�+?r��[�#/����x5Ҹ�y���o�H�lD��Č��V� `8���M�
+�ݼ0y�G�U�>��c]��s���W���u��Bė@�1_�f�S1	�������ѫ{-�-�,�a��M*�g�]�/��c	�0���ݳ$7{�H�4'3�tPQ���ai�Mr�0��/Mu`::\J��Bg��f+Ю{�t��_���$��G���O�'�(Jb��� ⯈�o7̎�ݠ�e���U^܃ �Z���L��9wI��xۂ�Db^�8~��"����
�pu��j;Sn�ctEr6T�c2!�Ct�s��S�O��k�Ќ�ߍ��ָ����R-�q/�DnCp��G(v]oi��.����6On;�W!Ua�����DL>6ss���h�s����)�km��Nit+}��\�Dm��w�Ri���ν[�&����x�*FU�t��g"ہ��˪j��`ƕ�x��K/zt�oe��Q%f1�t�jA�����걞`�s�X�Nu���^�զ�xH2pO�J|�S�,4b_="ǧ@F�K�a����%S��E�r��S���?��T�ʠ�\�:K����G�jg�!
K)��m�G�����3�U��z]*-��7@c7�	y'0�D�KK�����x��@�!q�<���w���a����8_x?����=ClJ5���f�[��m6��$�L�;+��>L2=U*�U�Ɍ]I-��LY�DwA�1��%�#8�)�kE��y&ºT먣 o�DԆ!@�,<З��;?s�M6�%�E���A��5��
�r U�����3�:$lƀB��@�S�׻�Z_|��g�¹�a�;�4~r�%\=%&[sАy�<>ϡ�����H�][jбmL���=��o�I����T��h��|�:#��4aM��ÀB�}�ׁ������5�����CQ
�� N2�U:.���R�O�R�����^ض�*��C��v�{�������6�)�ph������ J'�I<�{j�����%�Bk���~���~�.?x��=9I^76�[�R�t�vÇ����Zul��N�>�j�ħb�����0s6%Ŧ1L�A`HA�y0r�����L�*j2����`(�[ԧ�����n��3�:��A�[��;T�E� ���:�<z�CuM�!���?TRG�A�U|�Gฝ�O�PЊK@����#�L�Ѻ&i�.��9��3�8��Q�9�\��̞�?nR��/j␪�����! �]�9���zUi-�Yׁ09��zD��_6.Cf�Z&m:1���ɘ�D.2Kg�0�.�#�)[�:�M��J�0��#��5|aOd!�Ѡf���P8�`9J��3�E�"�d�b)֨�3н���[����#���5�<d�f+F��Q�	o��4���5��S���tG<�%�i VL��+>��*n�0��Ko�(ɕAB�11�ո�� ��SCE9�0���l���!���d�\`w�u&r*�#��k����9��Ӎ��y���M�D�A��S��x���z�+�G:S��UF �*nk���fP3-z�N�_Y��6n�	ǐ֛ޭʩ���$ڐ`��F��/\����F�Ǻ��Q�MIo!l���2m�祀�W��9�,+�-�2�,�;�$5]��p�~;��lC��WrE%6�g�<��s�o��6S��x���G
ؖ
��.�-xk�&_�i�<�h��1��G8#_D�kԠ�B^J=4T��$Q@��"�zv�|6pItF#��%�ɼ����*R? ���ܒ�*���-�r!����R�Q(�ZN��?�N��dX�����<1�4�$���oo8[W�T^{sb�#���3��{2w�m�ϳ�y�,����j�y�U7���A��w����<u)�<4��/�7A�R��<�ي��|���r䋐񐦛�+O4�5q����=��U�\FC�u����-GR���o7�ٵؙ#�O�T�D�N+��b\(V�j���A��$<��Y��/ҮL�E�t4�1~����g��.K�_��q
�TX[Z$�io����� h�Q�<�"P��ֵ��� Yh*�E{7�HQ���w���iy��yq��^���F2�k{�d)��H,%���d��A���.���P�cǿ��"G����3m[N)�x9f^�.R�8�>�K~���b�����}eǂ L-������6ùI-�����s�����Oq��4��;縢�ҘvTH	��o����ZK�)�ͯ�]�꧗�
C����҄gj�j PٞKb[�늍�f�~�+��W�^�f��.�XIk�'��ߤ�y����)u��"�{�\��GH���B8Sf~�t5��;�"� u��r��W6o�1N=Te�s������\����J�"fC-��3�hs=l���e�FEgD�c{N:�)�g*���`ee�t�|~E��g�΋%-03��C�c�O�`I�%��C�>�.Z�*��^�����	�D�1�SD�S+�+���B��ԕ�X;KW��dw���v?�=�P�t:�E0Y�SK��?-�l���X�A毬�:�v@�`�CNw ��z����(�������r�gug����c�Y줣Zܜ!R���7�|�==�NI��M�R� ����~niX�N��IBN�L��Ɇ|�aOUje��OK.��ʛ���@�$"Z�����Rˎf�g�&o�/5�$M��oSV�(U�����������G�yK�"����I���5�C��\3�O	�^�ŦL4V��T�$��#���2G��?���O6�Nf�(�K�>�h�X�i'��ہ2�K,��k`�(Y}S ?���>0F�l���=ʼg�V���1�=L�r(Ot!�y�MrH��������PN �͐f�ԛ�T�*7�h�|8ß�F+�ֆd[�ݛ�c.�bVg�]�<�;�v^,��l����
=����]f��rM*E\�����:��������*�Z�~c��LH
Xܐ׸����k�R�������Q&�W0o�~V?2���<���}L�b@+G��Q)�
"�� |5(�a&Fĉ��#@���FF���t�y�3<M-�U�6�9�` 	�uByI���&�A����)���9�'ƒ�O������n/p8l�aPq�9��vv��b��>f������+_K�$5�c3"��;h������!��^o�͞�:	�+�`W{�5��[:�Uv"�3>�	�㘁���P�M�
TP3���_Ԟ#%y�A��`��C�5l����.�� �7�uZ�����fj,�%a@�x��g|�W��	�Xn8ة)�zf���VC��1�g�5.�|U�2��G���Hn�������m�C[�j
Q�ѿ�ޮG5,N-�K�1H����o� 5�s����Z
 ��s�r���|e���ٵ-q1�(ry(}X-8�a_��$A�?��d�[ݪ�����b������˅{��-���o!�w��4���^����c��K���;�{W��`R���z}T��$�h�<U�͋c���*.gW~|�'���U���5� !l�Ҧ��:3��sW�����w#]�o�AUl���<�]㭅�y;O�*0�y��pj�D/���dY�h�C!��as����Ӡz��D� J�9����z��oN��w�e�o,���!��	�ǁ.I��|��U6̆����) �eZ0�rl�A�F#	W�dwC?�o��U�k<�G��D":Ѯ]�*��o�
��P}1M4�<��o�μS^���M�OR�e����3c�\Nc|�m" :��,{ إ!}�0����BP�+�MT�忣r}P1%�lJ�6E��Lh�V_��f��
�X��'E�Ή97�-r�U�.��\�.��_*�%:���osd�$n+���p>9i�q����y���bH��}�Or���l�l���6�:4������zw��kPv[*��N�Q�{�P=�u�
Pw9�qA�U�7����L��>Ğ}��E����z����vV��3�F6�I'y��譝w��ǅ���\��,�شũ��܌�jߎ���S� �� �����s��H�4	���t��V��IYi�.E���0�j-1���M��';�˄&�ї����V��	�۶7�[	�p�oҷ�|ݮm͂��:��A�X3`�?�:&�ȕ}߸a�"�l�s����(}���{J�]��˚�I*mp�F�Bx����4�B��d�E��!.�E��RVwHP�tJYE+���"$q�h_J4�T�q�u�A%�
����܃?&1�["1� 5��9p,�ݦ�HqU��F�̲o��M��a�Q�s"'����uJ��WB�i+i���P�,��?^�W��X�+�o��=��xu��M�sQ8��GD��0�}��lW���}�Fٽ�2�Z����F0��>����ӊ��]o� ˏ�B��
,-A[��Ѭ�~u�x����y1Zq#"R7��Q������|�jr�4����5��`&.��G�X[V'1�m1J�|=�E5۳���\��G %X��ڵvG��q�R
͕g��t<A9V�݀뾂6���0%��
"�:g�����6�ҩ��λ�8B!���<*ty�A5�&�Z��w��������Ւ0��D�+�
E�r�r�K�5�T�'Y6�$�<�K����/���V�d 76O����-�0�׆C�"߶����W����a�5
5���(���ݣz6��2��kn���0M���]S����o�R��)s�*�{��Bo�
��������4.�j-��0@m픘���'�Q$ �qA<�Z�v�
���#�@�q�?`z��`�HYOC�G�%��Z��x-Dg�z:�����LTQ"s�i�A���7��q�[�b�ه*�*�9��	�Jd�፴�!e"�X�µd��������9wP��'�R'������߸mF?�."�_��F�z`!9�TO�,%��w� 7�mn�BL:�J!�����Uoh�F0�{'�?e(Y§g���5��4��P��=�2l��e��m���G/���@�AN�S_)�.;2y�Yg��5L��6B�^���N���ޡ!+����a=�g��Y�� �"��ڡ�/��V� ��Il���e�&�+n5/<�N����9�*2c�wR�.�a�Y�W�����w��I4Y�� 
ArE����R4�J͙"�[���r��g��Q��
�n�CP�Y���0 ��0G Lͻژ�٫qgRB�Ͻ��FJ��ɢ)�� 36�΢@^�%x��ı��ʹ7 �*	m3G8��+$�d;�d�<��bEpr�ڂ�%�!��&�P��`������X�D]�� ��H�nvD8^o*ѵ�0U7=��0K<J��6����G���+�R�;
��s�F���M�	h�B�"�<J}��r�AI-y j;e�//�ƭt�m�A��a]�(	YS=���e[o�\�+�Z�l�ںNW�F���[�?� ���U��Z�I\ ��܂M�A�<�e���*��M('��J����Q���7� �Uq+t�	HQ�	�A�6�\������qRB�A}0Q���qkϫ*�3����p����8R&�5rD.QV-�l��f�,K 2�'�r�n�"���S�-͸.�Pȶ�~QFM��]��v7�)�ً�_ب���4Hc;ޝ��J0���r��������	������F�'��C{1H'�i1O�[�<�l.S�ˈ��-�Pƚ0���T�]�gfa#�'�էm�²�?볅�)�܌���ю78�O�o+J��
�J��ׁ8���~���T��.,)� ���Ӽ��V����fV�S����-r~ͺ�@�0�IR���Za�ଟ���$f�H��3G��$�g�4���2u�ʒ�51mǀW|��ؽi�������T
�+���������xv1f~�M�Q����`ؠ]��1><�Y�M5�ۼ ��!i��*�IE}��M3h������oR�[�ߨP��A� ����V�H.��$6��V�˖j)H��خ�q ���أP�����掱i�[�oP`��Ύ��o}��=��؟������l��3`���$G���_��cS�iI�r���0��]����S/����B9A(] c3��b�����˖���7��G'�(�W�$��h���_D��n�rn�8�E^t���Dl�!��[s	 �h1�[�$yQD���u��z���oSt�����󒾏�gqn(k~�%3�"�+lzf�n>\tb�aQ�y-5x�2�g�����;��9��aA	�^>�WJ��q��2�3�cA��v.8mI��q��A#�d�liܼUrUa}#��u/��r�;E�r@C��Dv�~_o��t�T��j��Yr'�5A�m�"�K�0�7g� D<��x4~�<]����p)x��fi��UIG��H���S?�'>E���}+��+MYu|<�<QK+!�㗶ɓ2�b��yl��K�8�u�ǔ@����l�^�a�'��EYE��1让��P\��p��ueN��{��R�������p�q¦�|=,�Т�Fp���̰�i(dY�<�JD{�,������;���[*� �����8��g�}))7��	�|9R8���հ�d[��� P��=Raf�EK̠�,�:�&ٮ2�	Ω&�L�tߔ���7|�;����R0,w7��q�Aۄ?>b)A�svi��6;���N�YKm���A��At�˿f��@o��F�-.�[KetX�i��U������F*��G�#�Cw-�����饫@L����vp�j~�!���������;��<{�;�g)Zק`�?N?T�z��C�m�u|�A��3:�N��bl�q$�ek8�����6�_��pc-��F�-�D���G�-N�:MgF$[�BQ��o��?�<M��-�}�F�����sw�J��N�cѱ=O-4v��0 ��'1B�R�XA�7}�4?Lwl��t�p�s�_﬍�~��m/��J��Ն���������u���lCp[��,��%�p��SX��/�D�鮺X�����}ˋ������(xq��A������v��&_K=�фEv��WB�Xʤ��h�r߾��Hƪ��/	�Ɠ�_A�^[ՄZ����2\N����l�%��L�⻶�?��mx�$�YtύTcDt��
����cUR�D������"{'�B��\��>��?6��]kܗ��;�9�R����-*?"sM,�,P}]�o��.{W�X�M�� �����S&��ʀ'��[ۙ��	C"W뽳Ƥ�$�thg��(�z��s�����qVM�Y����a��%% ���yꋙ��n�2A�91�%7;�����!�٤1C+��$��O�Q"�#LmU������,��M3%�%~@���4o�|�����9��D�]q�6�~&�ˑ��[̙���y�M�)n��Z���}3.ȇ�Q����	����l}����� ������ݻ�|	7ぅ+o�a-�@�
�3N�o��Ƨ�|)���"�!.�NG]NU�auK2��JUn�Ԏ����*7?8M��Ϣ �Q�8����������e����ٜ�2y*(;4L��r��U\��1�C��L���gi�7�����h�[)�&zK�S'��tG�q�H�� J�{)�
�d�ZϤ����Od�/�pF�0��OPZ_l�����i�t��� hO�UBh{u�x(r ��9�;�Ĕ}?�@�a����"-�1�!z�N�Aq;�_��N�$�����:�b�+�?�М������|��"��jԖ����`�V�c_�Ze���ˮw�Ʋ0�0��2K�n�e�;9�z�R}6J!o3����^��3Bl�y�{岘��/��c�A�Z;h|�U��<D)@]�����[ln8^��1zY� m�G~�X�`�]� �����պ�|bP�Q|Aj��0G��G	����SPo�+`�8���o*���k�����&2���%��b+,�ԗU�e��\��}�sq�#��ф;j{�=�!o)^�Y��g��4�[�D@ќ<��,/g]|B���m���	W�-%��G��Iƥj����U$ђ���Ϲ�!I�SI����E4��II#C��.@�c��ǭ��#gTse���"��\����_r<����Z��?<����d�^Q�ԨP�q��7]OՎ�.2�(VŎ	}DT�bh�ʟ������;ݥ��B%K�*�\1Em�G��\9 �*�/B���\n�p���-m��+L`����AW~#~)!9�m�{�Q�E���~
��}����VKA�,?��w��=��g`^H��TN�?�蹉�(NU�'�G�K�Fx��7�����blCg�J"�4�nk��tݺ��n�{�;,������sp�=�)I~���R:��և%���v$��t��R�R�gL:G��C�?I�Ws��Lq�4r��v��d�Lt�6C�3邈-�C��a#����J��Ϣ�t������n)YAq���A���!�Â��c/b��b�0'�d�;PI������E��k��ӫ�6�#�92���/�����W Q �(�b?'SW����J�94v���;L���J���� +_U�����ە�9u��9����$-�Xݰ�ky+��*��cb{��|�1�{����~��=�v��d�/��,�<��������^�U¢;l|[t�3?sf7'�q������۸1|F��~����'��,�����O���F,�y���(��(�ROD��)���j�#�j+��/eZ;��H~�d����]P�����Ď�ȺY��M�������vk��o��`^4�L�{��61�7v4���[������,�d8%�kμ���:kf�fD{��C3�*��sO�F?(�48�%p-���K�Aq�_���Yt��Ҹ9�;����`�͌e��~{[q���Q�u���*���u�.,"���Z���8(��֭�,�4�>2����<�k|9�q�~�e��[h�`}ݤ��%~�\�&j�a�֏I[i+�8߽}5����t9��,��yL�pҁG�݄F���-�¾�z����JӺ�w�\�K�����J�$�)����=� ��$E�"�i�M�	/{i�&2�<��Zl5�m-�":,���Y�IU����y-z��սќ�GKKDl��s�Gkˇ��>�}e;DtO/��jL��$������'���.ř 2�ؿ���ݽp�X��,�K�h��H�ٚs�E�PR��.���[S��x�N��~=z+2��a�8��SpH����w��j7K@��9.� ���qqڬ��Р��Hӎ���.�bS��Ԇ�\�r�̊ڠѮ������VTX΀��qS�^����#�b�����K��H��7c��9�(�ng��y\��|�U���L�Y:�,e���`"��Š����5��q�L��L�@��s48%���%R�]����-���c-|��Y즫���Bm��f	�A��,h6%-`�5��h�ٷ$�Z�R���L�|�w��W�FI�����%
1E�"]D�-�
F ��暉M�ʅhy�a�%��=Es��Q�f�%i/g�\ 1L�K�e����<<�#Sd�
��:c�'gT������K�����f!�$e`�sY�3��,I��Ys�t���߈�a:�OU�k�g�SX�q7��/v�l�ܤs�_�4]t�U$�y�u*����]-:Ǣ�q������u>�E#�p��=��������w(��̴A"4���)��=�^O��[Uo��b��X�y��/L����qi�E
ja�y���@��$�pԛ���y�9�;��x%�7ӴE�lO��:�H,�j��b ru^�����AP$�����b���li�u��-�X)����u�л"����1?Z��#>���ĉ��K�4�𘫝�}��E�7Y�a���rb�Ƙhm�\���h����؋��_���ʦ�JJ�� oϜ���{�8��	��	�[�)���"�F�x~M�
�u&7+�үn�V��=u挬&��������v�zyn��o�j5G���Qx|0jiw���%r�v$8��<���6��/"���|"l��C�Q87E�]M�B��D�Q�c�7�y�XK��O�J6U�X���v�y�DJ�����,��y�r�8m��v����3���$�1=.��A���ᒇ�35��Ў)~dW��M�6$��c���}H����T��r���k0s�Y�|�h8��j���;Ѝ@�D-V���G��r�x~9m`X<����4vK��__�Ȑ���=Xnw?�Zy�P?��ʖ�{b$�p}��F��uK��R8g�R_>bK� \�@%�B��vS��l#�j��|@w����H���� 
�Z��\������4�X�Fŋ,��Qm����0f���|�.Zj�9���k�x*�<�"��nx"#���r>"~*��<�q��"��ᠹ�Zp5��@��|�U�^g�ա�T_i7��^�u�Ych���ٮa����8�pG`V�3�o�>��d��\E��%҅��yzPl��j�n�D9թ@t,�]�+��4ID��B�Q�v��_N���H����R��Q�Ԇ���a������A�4�4��j�g�G�.p&�>m�h��w_m��-V&P��F�}])���#��7C�,R����h�V����r�������9�x���q���ӭ��3��zH����j'���f���F�ƴ����~����R���h
��#�|���v��]o�n�YS��A΀��H� �c���mI�$��)C��U׺zV�[T�V��$��tCG�x���F��I*);�D��|�߮�Y���9º�ōyv��N���� �w��q�����!���;�e*dT��[:_��k�d#*����:	6� ����פּ�Q��L����������旛�zg&����?�bpp�4`!'3��]�k�y�n��C��H��x�8>�8Ӷ�>���5�F DR|uV_	��k�=��2�}ӕ��C�:\�U�?�-NЃ���m�����Q4�G����6���ٯx�aP)��5��7��[T��3L�]��IA4�{�	Be����;N����0�F�G"�D_]�YB�*��@F}�4a��DV�	y�JX�<�^%�T�}��\|��!��}C;T/t���#N�m	����g��WT�(�I�}jE�����
a�#�U�a�`��d\yfѫx�,��$�*��:D�U�/�c&!��Z�*��w�{ ������yĜ��E���T����~1G�,�^r0r��I��4��b[�ޅYZ� ��3��;�b�E�,6�m��̙����z�H�C
^�S�A�ʎ*�u6�mس��C�F��Jً� �$V�t�p5+I��g��o��&H��\&��i�2�;��I���LY	nSD��w�n���0$������=�`����E�����~��1�VwB�o��S�cpc�iK��.qc�1[	��6Z{�g	��PO�$L�б��$�KB������r� ��Ř+�36r)a�&j�	��%��n[Yg�Wj�5ݧ[�4�:�q,[Ĉ�"ڜ=2c����wQ��,ew4[=B�(�
;z�a�K���9�������;�`��XT���w����X����
��?���YF����@���p�����S�|���+O����2`j��Iu�"�*u��X�\}LT�����=d1o���g��Zz���\L�Qxc�r��K����4#+����)m��n4C�$¾�[o�(�����l��J�K��g=�'/����S����tiú�di��*�HՒ�෻��l%��Gc�%-'�yz�K�(�V�1&fN���w��i8�d��U��)M��f�'$>���}���іa�k�> h��D�HY�u��I%f_�Kx\SW�j%hu�VN��C��2��Jwo`���lG������ʫ��� D<��F�d%+��vs��O�}
z���y���Nl�� �7e6�`i8�<��)%w��٩?H�B��_讑�H����'�d��x�
A}�Z�ԌZ���al���1Y��{����F��S/��`3�r/|Bz�f�q{���R��*�srKAUQ��Le�A������&ٖ�yh��G�;�u�c0/��1�%�h���+�T�s�ѝ�x��A��l)u�'r��
{q:�3is�m��Ԝ����LQ�WB��B��� �ns��r�+:I3]N����њ�"u��7ʹ:�|�Yŷ{Эb�1��E ] =]Ay��7lv)��2���(���:��khr9ZaDXO.���ё��
ʁ��d�o喓k�P��'}�(�&�� Xĸ��~��PP�;H�,��x�Mc���	3�jR�^��e��WZ5BoPy/HlR����y�r4y`'���| ����;d�A(Lv��~��1M���E�Ab?D�&�ܨ������$q�)i󽴴�.�'i8]��G�aJ7#�? �����V�v�N��P��Z;VW�Қ�I�v�E3\���bD�F��3*���x��G�8.�.���-�qJmE늇�뭾f��36B��9�~��&I0�+���; �����r/�B�1��_6��N���g�z�,\�+����f�z �OH�-.��c�y���%5��A:
����FJ����,�T����ș�R�p�;���/詯���M��hqI2p��������]s$�Ũ2����\
�4֍���*V�#ih�_��RM(��X�������R_i�d�@j)
�A�'�[�n��Qw�ߐ�v1�E� �� ��m����<�Y�@}�9���L�M�T�8Hu���M"�a[p�s��C	v	�}�D�m|��-��c��U�o������������*� �1��߇�ۼQ�}��%AƎ�z�l�+���C:����H����L���U�7��,�:u�Z�6?{b�2�N̫����r%������`�����l�tV'�w$\FE��[�Va:�3A�6�T��1͆	��q#�K�4������+B1>ש*Ec2� ��e�̠R._���[o����w����@�!׾ �����$	?G?��8����g#� ���+��7I�#0UۆF��[�6��3l��0�b���5Ґ<.,PD���t;�gz�^(;� ���M���5
Ts����2Lꬅ�+���?B)ڴ�+i�58�oiF2,.��V����y�+���A���u�������^�{�l)��祫�YU��wLd�m�h��+i���G����L��^���q!qR=��EK>]�ûJ�-��7�����-����Tp����*��GH�e]]�u��vRhH�bd�'�=����|^��D�p7�ny��"t��:>���U_b:�&y���^AH�ӼiPk�+hb~���#��S7&�&�5El� a���Y��2����k��[]��5�b�ʧ��Ӵ�<�|�l��	k��s�=��d}^�A"
��}�G�vO'���1��0=d�!��'���	�F¥دn]���%";�2W�ȟS�G�]�±.���@��y�[]ZR|ƬN�P�7��y����d��÷	T�A�W�&r��[ĩu���Z�2i"W��͉m�q�	�j|���I��[}BNn��=`*�����!4u#��P��C�k�sS[�m��Q�R��ͽ��MX�R�̐�8$Z��u�
Dz���Z���,�˅�J(SGD��q����cf��(C hpO����V`�euEȧdY��
u�=B�i����H���&|Ϡ׾�-�_N���8��d��fj���D��a��Q���O�3a�J��!��zmJPh����K�6<������G��zR�SdD��vm���C/`*�`�\�z��Iʟ~��~�N�{����+�`֕�~� J��rdU\	rf�WP��ň��7���6�q�{3X��7�����G(,�c=���I��@gOf6�'"P�V�xr���u,,�/� !�\��+bq��w�#��z��i�`ͶGj���b��� �.\	>����Ώ�Wh[C�6�*g{�'km�:�}9T�?�Ə$��!����l�r9g7[�od?I���m4�"�lA�NP��������?Q��U��X�!v��+�Nu u�"o�-��� ��3m5} I'r�8Y��CED���Ab6!p�W��w��	oj�M�6)A��b��g�p@��m���E��e{��^sV�Do�\Ȉ�-"M���0A	]VGgqzՠ����Ph�D�Uf;U9�w/�+�F�&��
�y�Քר���d��#�@����B֮�'��S�G�zذ-xP����������2x`l�iE	�:Rm��ꫨ�!,\���v@78ևp���/�qp��.B�D�jXtW�w���H�k�0���&z�+���Cl����J�c9xp2KL�'!�>���e�����g�D�Bky�FrY<�Ϩ� �YA���yՃ��$����=G�Z�j���"	��_VDFcN��#O�bG�3s��H�������p3��?nb���e��f�N�2;�ʶ��c�)��Z6ܦaPR|i��Y���
��-uc<�=�k���֚�oCuy�^����.u	�|�m�7�36�3�O�.��U�^���M�7U�9��ig����VmHHG���/��~a����Фd�_=�U^��iB�>�K�"�c[�Yb���yQ_�e@OM���,c�1'�V#I�6D��C��y��:^��{���ơ�4��&�<@�%��qY�6B�'b�Ãe��z��� g��x�X���)�"�[D�&��K<V��̑�T���j�%�02ڮ�^��d������Q�U�5A�,Ѫ�*��V��LMe�1Ḋ���(���>�=�vJ2C,Bt�H�,��d�Y(0��i�;IV��V'��Vد���`����(+�<e���x��IAyf�B�}����
�{�"��`Ct��))�N䔃N�$K��Cj�p`�O��2��\,~Q�]�"r�q�T��Y�B�PIT"��{�L�ə܁��E/��J���R��=���v�Cg�|)�3<�L��r�ݮn��Us{�����	��T�e
E;f:��LH'G�1�'��:Ջ<J��nQ"\7.�v�m���*����ظ+>�*�/�m)��y�����S�Y,b&��MY��u�&?ʕ�-�LtX
��QR����ރHj��~w)Jsk���4Y�ŃF�W�7V�<)jF�\���D�ct�
����YW��]�E.��R�����j,��6j�Tb9�!U�[��)�FO�˿�A�����Ug�^�37]��ϖ��L�� ���κm�ZY�����Y�Fy6�:�r�$�U&	/�7�)t5��!	Cz��� �pʅ��MWB�H@��D�`"�N�r��Z$�������{�������g��Ab��i�v^�����E���`~��Z�$KD�Û�Ǝ�'٩ǂ���۽�����p��ѵA�f�� �C|�ѥ�˿c/�.���"D(�H<��(�w� W�G��L��Xlz�ߐ��L��4����֭��T��ρI� �;��p��&޵3�o��^�&�R��6�v��f(8�T�����w�$�X㌆��sā�`c�r��Oa�J��	�~��N+��JZs�@
��!�W�-'���<���H8Ez����7� �4����d�WY�2�]�l6����]��)#��t�VE�� ��#}�]{�e����HQzZ�jКN�����bp�q�FX�Aj����Ѧ<K��^���Tv%��պ�F�`r8
�?��D�9�vڵm��o�,p
�zg�
������H�J��
BZ�\���Iv�C|�d`8U�Οi@U8�5�m=��I �&��&����C±:�醌�_z�1H��F��m�;�i��J�5��'�@l[�	��<�A!��1����m��,��4�l��������X���'�gYa��@����(�<R���������:~>����M��Z���o�G�m'`���/Fr�V��H�������_�����D��!0ec�D1�D>���~�.U���_�(fC
��SL����_���w���D(�{�wn��z�W�{�% ���t�R �kH�/؋L6��f�Y��]_��G�J;:�I��Ż���9�7��N5K�:捒����11�U�1Y����	w��h�Y�	V��t
�����<����=����u�� 0�,��H����K�Z�4�Uɮ�ށGs���᭧j�=�k�zO������A:d���aIˣs��d,5ևG���ଝ����Y~s�ށ�!A�GD�����P�T��A��>����g�t�~�	���Q��`�@�9��D���O���xu\#(�S�܄���EiM	H�w�k�_?|t����E���d�|r�c��C��