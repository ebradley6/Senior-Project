��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d��p89��N������Dacf�o��!$��Y���*�#�`b�[2������T��Y�c��iN�7��3hnc��j��J��c�ޤ��������t*���a�G�/���1�X��S���0R=���]9U�N���
�ݖ��� ���������p,��F�Gb	 ���5��G��r>��T�CFQ7hQ�fr�|��H9^(�K�L��5�_w��O�R���ƃ\)����t~Gf�;�x���<R4�O�槑s8X�z.��DC���o؅�>��,f�n��4����-��#hp�&�1�*�.%>1��"�hn�@��I��yq�s���9a���L��)�����2d��� �tpi?<Y�������'t �a]cn!�-�� k�;�O3o��Nܧҽo)�J��"�m<�u<��iB]N��1�{� ���ɉ�P��D�Wl6_�8��$a��%'
���'U�������r�[C4��w��x�gZ`�uZ���8!:�N�"���%6oN�0��y�Vd�Q�7�-�bvy��ގ��P��!!2��_U�6����A�q�MfF�j)��`$��ٹ Gd�)e/4�(s����$;�Z�R����f-l �M
M��]��5Q���Pf�ת	Q�XK�x��b��}�K>ח�5"�?I�����Uh����T)>��2�(a�M��`T��˅$���OpTH��������39�S$��E�i9n�yG�	���喘��_��@q��B���@`|1���>KD����kr+���C�{�i�R,�mL�
M=y�����>��h:7�ż�������N��R�#��-��?�#�Y�+�� ^�@�.�ĥv����'�u\{��d��Į�&���8��v�Do�0��r3]G��Ǳ��\����[o���@�nD}�uRa�u�]v쵛SK�'<戮6����-�u��6,�F��#�0�'�k��O���a5q�1$%��1�� �z�c�R�_!�m��ǛK$�O��D�.���l?-LKw����E�*��>f�`��:]	r� �u,�R	&*�O���n�DE|��d�K�s5S��+�)."��N�g�L��Ҵѯ�N^�6�x>�/����(h�u���>b����i"5�l��� �l����a,v����\}���b0.��=��1́2vG?Z��o�\r��H�IV>으o���#�5�\��
Ʉ�D��E�m`P����u� �|�Ѩ0o/�Sy�O��x���ü�� <�Mj�C����=��"�FsDz0�22ZG� nǨ�E�&�&LbE�[��e��ƞ9��8��r�燫L�l���h�C@��X�'CV�x��L�+�������P��z��p��q�/���*�����N��'���p���|�*�L�t���V\�t8Pڛ�3
�S?b��ՃSg<r�þ���\ab�No�U�h�A��r�Z������+l^�^������sW[u9Fm�'OB�[�7��v>�"M�E)��Se"=�f(�|e��3�-/K�?��NJc���F�f�IRƈ�u5g���^Y��J��ym&9Ȕ���Cl���z\�
�J�����kB#��4��~��2�+�v�E�_�o��sU[�gg��R�������3`E��c>R���~�Bm�{\�/��rj�D0Y~+��?T�UCօǚ�<����+j񵇡p�������E�rс�f�<Z?����%/#����*5)v��B��X���
�m�T,f�ם�\v`��L���C�P�����qrh<��8�A�J�R����dR�ԏ���yK�es�u���^yu�a�^�:$�>��/�����q>?�A�^�)������ޙ�+8`x�%��ya��z��Ku,��}.-`�]UnB������cW�B'�����UT��Z�|̘��~i.	
��������O��m.��$�3���\��*�~�7
 �#{j���uȸjʐ���
�Uϸ�]�T�� ><�@s�6�u�R"m �h�*�|��5�N>42��;��y���L�v��|	�4}��zQ��3)�-�j+ϑsT��[�'����l��J�����G
[�wt<��% �����v���jL�{�`Z�\p���0��Nlm2����ԦN�I��_��tq�ftwH��QȂ_��$K-�g�B,R��zG�A���6i�Ú����B�ɉ��"��-:'h˧����y��'���r��HF|@d$i�!��=�ّ�^�[�"��yΓx{T׹b��D� ��4�.sD{�S.MY24���ԓN�B):~[U����g2Ğ<���K�)�-�a6!t�T8���\e3(�Q�9�E�!�$��u����"��/��߾�f���k�R+}����~�
 쇒��\n:�%�VN Y�fVl3�ņ�BИ���'�����v���:ɎDZ��B�&�������Cd�D��-�y����6�:#Cr�毟�a72_y�"O P8�N��^�#�:�ҝ}�|>���?�>//� �$|���6Tk�U���@D��)�����A�-ٶ���_��BpM�	f����.�w����g�]t�0��|�Q�NF�d�^Z�s�V]�JE�,Y�����`_L �}����HQ�%+9u ���A�T���ܱ�Xa�VO�I>>�mTL5 � ,������ٵ$�޵�ZW׬Y��$Ca���7<|���s��2̒���_�Uq�#reT#�V�E`�L����T���M�e���N`M�J����&����l}�1��U�@�{{2��D�i(3ϣ���"�1�I%>�@E��,+���r�s�����֔����;�¦�=�%CBPo���)E�R�S�..W��0��d��$������p!3�i�zG�)�q}g�����ҥv�%�Y'��D*"��@���kj�0��#m�.߄�	f�g2�oc��8�8%5�%H`���1��LB��qDgt7���g��-�\(.������{h�Z^�n�좖�@�ڷ��q������E��8F��X��ֺh"�n�҉9����eC�$m�R�u�򫼞�d���hR2���[�
�6�����q	���Ȟw��~�G��&���z�#�4�2@n4���7'a���(!��5�B$���(����Qp9Iuv3��R+�l����q�%m�̹�'$s���G�NZcX�CX;��Y©��Ut6H����{�$�@g��L��*����G�Bg�\�f*�e�/D"G�vZX�7F��a��N~VL u4ٖ�Bq(�e���y:�������rԣ�K����`y�JZo�B�N���w����2�Rl�~9ֶ�)�lC�������\G���Y�������|&��tY�E��x4����U���+QW��0��پ�����!�o���-qE���I-R��@����W�-��^/o+uA/ܠ�����б�ɜ�����|���+"�:���C�i�z���bK�z䵬���M�[��� �[�r�i��`���S{|���*�8ȱR��>Ys4Vd��L/F�ר
�B�HDQ]`�q�+G�~���>ki���Ss�m̠�E�Bd�cNg{��g�	��A�ǭD:7~���W���Eiv��]�i����8S�J�3YZ�l�ϋ>�(��{�zÞb��gn���M��E��c��|`SXZ��WZ��ު�d!��Kn8�	��<��k^�L����ҵ�!�����`��$�ϯ������e���@�-���� �@�n��1��Ï%�H��j)=�`��{n�Y�4��΁�\8���v(w�c<7��Z�+�hE���5�#�515(��G.4U��z����f��`o/�Ҥ��8؉�N�{��t�V�,;�"��g�CF��/U���	t8�H3EM�����I �I�j���<L'f"�]�� ��f�i�2�%�&�1$$u��T-m�p!�����ȱ5�~#D����p��0�CT����Φ�휠y��T{���������ÞM�PF	�Q`xo���/ ��%�fusMs���L���d�JEL9a[���o��id�&%��l鬻@Y	ĝ�Rwu9t���v����|����̟�?]�[3^������f���b-�W�1��k��cn��b���?�##%�a�.�Wx�XU���]����'��ތ8�S��5�	�#p�{���]�%��(
���f_��Pȳ�qP��8�����6ԝ ��W�J�p�	���-H�٥�$jx�$8<r��6
Tgd�v7/}�h'P�n籘���+ ���;�[����[���C"�"{�����M�ѭ�a{� ��U�y�[=}�&ҙ�*W�jF��fA�苬����I�/��Y���b_l�F�_�u��JY]j�a�>��K��+]f�D�=�=�&�x�w�ʩ������p=, #>K�^^$��� ���+��^&���qT�zגs3}Xi�E���!;����[�ג��a��U�����ƥ����jޱIm�}uH�5�CYLF��u�1��j �ֺ���zw���<.�����,s�d��vpq��,�����G�_x֏S�c8�Ai5�ɘ*>�����Ba��(a�ie֌�& �?�m�%){�
�#8���껽P�/Q�Hţ�׋�`G�mrN�� ��jyeM��� FX�:rS>i���w��e��u�BP!^ ��_k��w����r��DF�na6�T�Y��X}(���#�l�$@$��C���q'Sr<$�- �iU#�&�����f�Z����uj�xM�;��F,i��� �Ч��<�0��#a�68B�DP�f��M�r1!^4�Z ��m!�!_Y��X�*����L]t�����S+  �G�%`��Ttg�	}�?0
��I�u��� ���C13�#g�*�U��}��OgIs�HC�Y�ځ�_(�����5rӡ��0��$�~�)@���{��)FL懢'�D5�vI���S \ 6��_N`�
҉@ӄ���g�����V�j�:wfB�t� QQ����BC����8�z����#"��26�УtP̔{�Y���t4u�M��>��[�%��>ƈ�Pm��M–��,��CÓ�w���wZ�gT?�TmЖ��D�v"��W�������@QAv�v�u'K	��L$�ٷ{�b1��4�!\�Y���Й9V(�q������N N��fC*�����\����E?�E��"���z���B� �{U�y���/
�sp��ݶ��D/p$��&^H�]ǫ���B��ġg�p]�@k^�fmӷ�b�S� �(��-N?+]`D��)9[�+j��]� ŭ�CC���:�<�~i5v�Ӄ��x��-M�	����5Riqu�|��eR�I'	;��>pk*�<FZ@͡��|�[r���YDoa�I��C�i�Nw��.����1�+�b�Vh�ZNc�{f��]��>c�'�*����U���\�0���W�N+��Y'�U�F5��v��}��p��i;�m�IG�܋�#�a�̵�i�~Y(��?3<l��-6*^QA����y�j�jE�~fL
����A��s��P���&OW�P���o�F;�/zY����y����;�!�w��mSW�i�rh�%���i&�1 �ʽ�/
*�"I�2"\&O�^��[Pq�W���[Fx � h�9��vƕ��_R׳X���:��P*[=�|"Eiy{F�\�UIV�������8���W��{�QA�ہb����b����������n�y�Wl:���/���U:�k���ߘ]�n�G�@[�#�^ ţ�	C0�L���UO|���)�:o �}~M|�3�j#�A57��F�W}����.�̵�*����[o�v�<����Ǩ��E�h�Z�@�?�AN�R���[k�f��\���+�����oMIH�Ȼ;�k�O��ϤC��c�Hj��U"��[:Df�n�A&�q�.Ql�C,�7̃c��?V��e3B���.*4�m�xWt٦� �Ę�'�����]��l�g��=l�Q��,�6_���B��߮��@��3u'�P�o�|9qW�;.R���P!��׌i����`� ²��Р}���yTp/ۃ�o0������d�5F���_�w�����˺�)��[�A�P����q�'C:����yH-JB�XJ�E�A�`�؞����(}�+e5g�"�����"}��-�ga�(MFJ	D/7�J��&���?Řy{<�+��V�/����F���Űח�!-�k8.8�j�q���yMk�Y��5w��]�a�����i� c)�Z��N�N��Fx�,��}�i0v� �T���-�[�?��r��㞵RV��rkKn��F�r$�(�����q!�_�A��7�5@���� ��'���D�{�[xE��x-5U^����Tjի�b������إ�Ѷ0�b(l�y+�e.�����<K��TI$�Uxa�����\�+�uh%FՄB�����/4n�^��:T�[=�NA�oT�R|�FF�kwr���K��� �O�����9]�C�R��0��_���(3Cb4�
ˀ3I�M`�w�`�B���ˈ"��/d�+�� Jk&C��>����ӱ|��u=O�G�Va����IG�=�.jZ���Q���d����n���{������N��^���]���v�r7���b6l'Z@���,Gp��X��:ѱ�`���ց�����:����R�4r姰W$�e��"'f����R�y-�ۏ�H�T-�]]ڸNA�e��ʻN(��C��iw"�)G�	:�7f"{�~�i�@�/.��|��2���oe�L�h���˾�$�z�ae-<1TKu�z�ڽL��?����&G����p67��&�0�.��ز���{�P�#��si�?��P磷3���TSt�_D������}��$�[<C��nq��P9�\2��VKG0���܋�+�>��Zf�1� ��,���h�����ΛP���� �+��t]�!���hz�H-�r��5�Y�U	��*b�2�,����8i��B��̋�Q��?a����0��+2�}�#��n�Xġ��;8��4�=�X>4f%��r\�c�J��=(g��ѷ3�?b����M���_��C�?˽�e!�(��D�do��	��e�%�#N�"���hǥ������a�!��9��HX���1�D�̌8+�Jq�k��X��`]��0=;7]ե~;�"#�KW7Y&�P�Fr��)�?m]2������E/���u�52��ˋ;�N��n�\V�I�����Utʃ���BM-P�[�23C�I���V>`��s�x�&h7}G���,^��%�^�MrL5�זZ�"h�����Ѷi=~��9;q�Y��f����j�ˮ~��<�1������"����	f�(����s���}��8�a���a)4� �VWrS���&����o�c�&W�e�UEP�M�B��K@�e�2�4JLsaO�e��q$�͝C__S�������c�dFT� �CnCGK�	q:���9qȃ�AgN9$3I�~���ӡg,�8�7��mԎb�2��.o�[���1�&�\?3�'!&����]�y�0�a�P��[��	ͦ�A��I�~4�4�pd�<��q�lI�{��u89����o�Rd�L�^�fIr�)�*A��[r_^�!�9~=H!ΐ�A���eJ9-�At���o�6�{�6�-�B��ꞩ��R�M. ���o7wfX�Q�xi�%��S��ac�[2��ҡ��ܴ�;ۆ-r'�DA���|(C��i/�y� ��FJ#u�=���2a�Q�|r��pU4o���G9g-�<�B�7��Rh�<jy3jef2l���'	)��A����Y�סȉ���8>�t�����<n$�P�q% �(����iw��~f�/9�K(-f{�A��I/ҜF�<��&�u����'����=�,��'��2%zu>����[�n���<\'���M�� {<J�m}m!(y�{��5��%�[�T�|�����-�x@Յ�P��	n���)#c�~ z���$�A�B����gM;Y0�}���#��e#_�cZ��Pt�_���v��s�ٶ֪���	.~H��{F��#��� IAdA��M27QK5�4��;ٯ�\q�yR�Ȥt�p�;����J����b��Y�=!�Xf�Q�=�v]�?PX����2�@��
�s��Sw��JS/ 07���g�^���~��9W`��=��=P5Y��~�����L�=Sv+1�Zs�6F�¡�Ҷ�,�yeN{�����t�8���{Nws�wȫ����A�6�WI;��0��l���� �Tk	$�{!r=⪼�2e�ˠ�"����H���ŭ`�@�T��-G���.�5F��mOQ]_VsB@p��0��`h�o'/wJ�'� �s+�P�^"4v��1�RZXj��z �>&�mb�Aߘ���k�VYV,���@�/8�OoC�$XuD?kN'g6�L���H��g����n��RD<6�Ӆ�c����[����9�D*��_�H�v���b��:��m'q߁ �-�O��Nhi��A�Z|@�ᨳ��{;��@^��0�&ؘAa={Ӯ���i<�N0P �uk;��:/T5ʲ��_g��J�:�aL��B�c�¹Q1�>�_�/��F�"~��Iz��8��T�i80HK^�Q&��ֱ��[�d��E��Gh�P��YX0_*uW��E��ƫ���N]���0n������z�Z��RPOz����N�Ҙ��������c�
���I����b��񰫙dpS�)�]�����Qs�2k(�qsw�crq����I/r�͞����\S��n�Kg�8��7�+Q��"~
��*\�� ��jJQ���V�{�KDD�r��VlI�i"a�,=�f"hcG2d���ё*�d)��Xl�(FVmY�=�D�g$��f���ե�Om�`��2GWI�=��4(`�v��\��y:�RXIü��y*�\a�ZW��_U�������� (1��֨�F��5�@�v�!��H��Zέ��=P�ܹ��NH�(�]���sg	gm���-L�A�1ݧ	��IӀmh/@9�Hݦ�[56{5�d̔�w=v����R-�9`=0�St����zE^0��)�JT8Ќ�?N��y��H�t����y�5q��r$8��Ck�N�{
���`1g˖��t:����6�Y�����w���9�ދؿ���V�y������Yr%0�K%M3��\|�U�"��16�;�.�<D�/�fMu�Y�s_C���gz���Yu!��N�����a�R�HJ-�A��'t�Ck�\�8���ñ��"��{d^(�^����#�0���(�B�]ǃ�`ooIov�7���8�^�����VW�[o�$v����"`{JQE�h��)�5��Wعr0%��r� �W��	(-��E6�T��/�A/i� ˤ;_���q*H���fλ��?�h�9�z����ǚq�7��Q;� ��-��̼@ �L  �A��GZ"2��Pr�)�Ū{���{I{r�	�A���&w�>ݺk}���iNW�GQ�^�g�[&������U�^B�8�j��)@<�Ud�G�����e����c�E*�V�T}�}�N��ͯYٳG�^��N��Õ'�n3m�2�v�z��O����p4�����Dׂ/G�����C��R�Ñh-?�e@"-B�!\��>�c�Q^��_Lq���ڽ��K�� P�*ص�6 R>r��B�6���9`���*�:^!��z�O_����� �����x�q�x�n%�0��IL� �g�$���A��������P�
>� �-l�%~�������T�H-<ӛv�����>��2��7� �3�i��:T0���]\�$&W��d�o�y|���v��l�pM�;�_�LX��&T.�����Đ���j�7�Qp�Ŕ�4$��s)48�3.��e�ȚӬ��L�)����������&i}�S���,� ���P$p��$�˂�'1˧��o�oMD�B��]��B<�$��j('?"�IPn�l�y�i�}y�oRD�(��z�2..�?8n�1�[�Zsd��ك@_ez<����#!�����S�%�����\�@ǜ=��Bcui驩ˮG6+�`~e�q���A�&r��J�W[�ݽ�w���+�lUn�*��cF��Pp��B�U�S}y��J����p�H?O�K������L�8�����������vV��{����zTG5D��R˃��.��'�] �-�\�#K����LFD�$Q�"?��)o2��
�;��NB�x��ߕ�6я4����uA��3��qԖ���w?��um���{XS�,/�57�5^W_*z�$$\�<7��D*�Y��,���?H]�쌮8��e��H�2T�$ꯂ�dlG���_��Lאi"����OtQF4u�j숭v3Brj+�
Įg�-�Z��y�@^(��ر��B�͘w������rTI��"��?���񥿋��xY`�ə�x{��꾔�}�kS�|����q�S7����N���Ah�W�}���>gCN-���C}��#kT9=B�"�"wF�n���J���]*p��$�4:JX�jwO6enU��)L,<�/(�K��|�m�wG�}_��%� k�L`�
kf�u��Kģ^�_P��Q���K*I_�7�*�����Zf�S�O=�M<���v1�lI��_�ੲ�%�Vg�ċז�B�hك˃�['Y��&{`�<0	c�瀹���o��FpG������?ڡ�*�27y%�E�K]Q"�>f����[��G�0�+���ަ�y�H��=&/�1G3:��� �  Ч�{���W0���#����æ��դ�v��y@<F�&5R��4mò��"B����\�ym
[��tH?�t�{fd�)4��e���v�\F4�H�:��lA�(�v�:/�w�^�����S0vXq� %
�{�9�"�V�%y6v��M5�%̃b������S��(p���b�4�jM�&�,!eS�=8��wX�9��K<��-��U�9���4L�NE��k�	4/�]OҎ� 0$t��C�����/I�����σ�Ux"�EH�'y��)�X|t� l�^i��G�0>xn�ݛ�B�7���n�9��J�R������VH$��L4���N�7�w��dI��O%��I�>5!��KwEF�Ft��2���e�.�)�����qa��T؃fX&����p��Bbr�m�D�8m��YW��L4V� �4���7�(����Skg�@�
�C�E��O�칎�[UcU ����f?�TW�[v��O�V�I�JF�F�b�4d ��H���|���f�Ld��tud�w�β;5�����!��|V�X�ٹ�tA�Ɣ��%�J�ÑaQ\\7�Yօ�6�@?�JT��f���WC���jG�f�h�G��ݟ_5U��#q��[���r��j��u�.̉���@�&=��+j����z�[�������q7��N�%�3t�5�n�=uݶ��z�y���3ZvFA�pBu�.�6T[����WW��!P����So�4���+j'����Ь����'�-�m_{�4��ԃ*B��C�ZP$4�D}�I���o�D�̯���2��z5�h�yj�QQ��TP�[YÈ�/̏���Y����Pe	PoPȆ##V�(�o��wI(�{�y��LL��%Y{�CͲ��߄�o�jCϜ�nhX�u���P�H/��r,H��bj�
.�ђ��B��N>�q��������W�@�$Zd2����Z#}x%�<��w���4������[wJ�V�%L���۔���'g��]�2����@A���F:T毣]!A��s�J'E��^�И�Ғ��%����_�Q4���O�5��H�:���̔z�S���N��/ ����#�ʯc8-'�a��HE�4���\�q{�~�p��iJ�� ����X����tD[� �F��8a��MR�ћ��N�@y�9��B5�#1� y��n
�i��cS�Smd��/�цg�z��pf��j���H4ӈ�ߙ�M��Ӟ��B��-ۮy��ѕ6cA���洩=ȝ�`�=-��S�P�k�qZ׎�r�%*�\�<����3�e�+�&���sr+�ֵ���ئ[�y�d�6�.Q�`p����<9h+����}�3X�/CEuYB�q���R�o�HIWiI���L?��r�šD �����^o��$6c!W�o�B�04�b����R�,��4K�I�{k�0B޺���-��h	��� y��,Vӄn���<�m3����I�d�ܿ>u+Sǿy���ޒ�E�g��N� X6��s�<C����L�⵾e��|k�h�r���@��S�;��-B�n�g�OC�����.����:a���d�%�ӋY
�W�
\ϣ�0v`3^�"m�J�P�&��7Ly�՜�3Ս"��16�;�
�w���+�$�K�,?�C�D�AOv#@c���UY�7S!"�9����9��]_ȴ���LjH�!���� ��T�N�v��sV��eb�@�r/�(�߹Z��-�}�)�}��V�D��6O�����Mv���o!U���RMT����P�1SKfzD�)�OBC*�3P���$��L����XD3�0gIFb����&�`�:���<����, ���E�"%��2]���^�h��<�]4M��o-�,���Eͳvt�+�omr�e��7V���Wj���I�zz��;k9��[@UX�xЍ��W-e�U�����iԉ�Eg�C~��|/j  g�!r$��2r���N�*���0��(f�4d�aE�Dc�>���ef�WmY��6�����B�b)1�7]�F]��Y�_����M�W}~�+�gS�C�;��	�+p}�
.��$��A��ohڒC<��Q���ve�ʤ�(��G��1��
۷��<Ҫ�|q�D�W+@,p�o-4��C|�P't��Z��_g:�4 o�U���U ��Y&���cӌף�@��9�$�Y٧�۽F�������H8kRl�L�LGLŻu��sE�4}�������%
�#OHG�s��e��E��#K�e��RK.�m�=��^����4(����Ji��(|�� @�)���ZF9j�+�?h�'���`�����K�%��^��<M�z��D���Z2Q�72j��E�'�Rd,����7G=VFl�څ<M�#�5���8ã�x�f�JDz��t�
|��!��G%JgX�
ȳ��F}�UJ����Әg*p��?3������s��������% n�+w<M;�sb�^m��	$�6�������D��?�c�AS�SmO���9$���G��a1���pe����aKm���w�r�O>�`�@m�
�)*�1��w���7���Sx��B���"�~�)8ր� m���>U���2���l[�ya|H���Q��^��S��d�r�,8�p~��{���qW*]�
�����-G)��ϩ�=�K�}>�U��=�T��W�Ah1��D��0?QK�8��JQKu2��
�ĽN�J�0��Ce��A��u~|�d>�9�M���7�?�3+ݞߕ��(�]�|�����[�y�Oփ���G�>���U%�4�d��qΏG��uP,�˕���l�n�d�Vp��64+N�Z���p��'��m-J�$԰������9�0{dt��x�s�P�D��JZq=��8Q�z��i3ĵ`4ҟ�y�MO(�{кJ)�c��?:&M�f�mET-I��睳xF|"B0�ՏCO�^=XY ��E���麶/9Bq%���S��]�`��5_��{��d�@�����ǣL'e��zy�(|��`q�����\B܄��86 ��o���u��R�k9Y-�|h�?U%����ӿ��KjrPnQ�E�te��>p�EȐ��}���d�%���8�č�L�c&��sĨ%A09��bv���qx�U�ƟC9@F��������ܹ}�Fl&���F��=mR �-�mk^g�vλLo�J�K�.5�I]������c���y�---wl�n����)K��Qq-�[�ɆC��۵^�A�`�lD�ג�x"\Мo�6��$9�L�������i�"��1�u�N���0֫o�S*g~�Ӧ)�$U={c����}��������͒�����]>f�i�@�&]��z��:��i 翃����}8�?5�r�,�3��_�>�j��!<�R���B�� ?K�?Gw�=���mt��BN��v�)�C�$/sq&�
�fWL8LwaKg�_I����%"M���%Ef�(T�c��Ku@/KA� ��.�%�R���3���`�޶������^��^;�{�:yd��%�G3��)� �vk/2�%ߚ�;��_A-m������Ϯ�#�9[���S��
X|�M�ҹ*5��lywVc#�0Z���[��M��1��0̩���ױ9��ĽR��kd��A����QP��	 u5���M2�A#��-��4j;�Z���zd��O%Tt��a��#Hd�����۩�N���E�T+0���mE5L)�=�x�lUYM�؀�y`)u6�˗L~2|-�.H�<ʎ���n}]cO��ކ�ڵ"Z�������B��D�-n���lTT�-̀A7�����Ȁ�46 ��KW�+s|%��e?^dY�ɑ>ʱ��Q���h�eZW��쐕n87)����T=����D0�L	tԱ}wF�'���H�2�].a�e�b|�ۄ�MH�0Q�i�0k_�r!��Š7f	�|�:�N����C�	i��� ������d,B���\��o�b�~P����:��܋Kոu�EiY�-��Xnt�HL=�i��|9=��ɦ��]
�}�8�X��V���%��!H��2��]�5V(�)H,��e)U�����đa��"z:�2Sk�4(�[u�z���}����@�������s�x��k�l�<���z�&�^���dtI��a'ROz؉�͢"��Lྲi�\��S����>o ��E�_Y� 1�3���d|��]h�)Q���f��sb��zX�^7���Cܼ,~�,J+�DĎ��!�� ��	����셣0
����$k����Ɨl���}3�'�b��V�L�%�즀ܷ�7��$;�3?�e	k1*?�%57��S�P���K�s�;p���
�e���d\®��|%�b��v�i&)<�g���5��l>��W3��(��r��C�>x��FS���<�����!%=>r�
���wi��R��aʘ�~��h�����.n�!k�d��X��]�߉�q�:�k�84�M\f8�a%�TT���n�8GGw&��ez䅩��o%��Q��q ~Zf�9��n�C@��a��Z��I�vg���i��W%Q�hZ+�6:i��|ӄp�;-�|)��`���M��J��!�/��PA1��C_�h��n������2t���̙�؃N�Sf� P��6W?���_8Y�-��6lN��t@�#oy_CL<m���_ȵ��d ��XQ�5�(�Z���gJ�g\��h�7qZES	�Ď��:�b�P�T��C2Gy^9Ψ�����2i��y��sg��˞�o��B��R�TI�n3���_uZ�:a���U{C���T~6�A+��K��y��Jz����������ീ��[��j�Gq�=��h�����{r���L,E=��� &+�����¶���%��<̘�}}��*_|��$����T9��j� Ѹ��oX���=��(ԫ<϶���+O2��|t��1� |��F���������`9y�ġҠ��P�l/�,�p�r6��έ�-d��s�9��OI�����b~{a �� ����ƾn���f̲{7����ȅ�y"�"�eWa�FL�~���*6)�Y�}�mr#h5u8/��jZ���h\	�6��d��"{Q쑕Hmp)��u��p+����g�Nj0T�b�쉬��|{am���D��Kw���)r�!
%��ʞ�lHȘ��%j�T�*54p�V�z���K5�/}uaQ�S�D�5"����� ?1�ȩ�4E����\�*g1���UI��ȫ�T��^}��-Eu�Y�9�U���@ŬdO�l�>L�89!(��/���D�ZMGU���PZvH5��_p�-`w9��
�)ps�q��:��7d(��_e�W=�R�����4UaM��G��$Ӯmm���牦Oz-8�q����ta����̀��>�wZ\��a�p~��ri�`������{V������Ò��)�i*��!�k����JJ�ĮD?�O�K�мT�Y=FY�wB_M�$HO��x�V�F��! �:�b�^�������D��2�� i����3Hn���3��)d�i,#�s��w��Z7�!պ�Y�efkZ�?�ˣ��偱q�FA|**��c9�L8��Ft8����&��X��6B�4�sy �˞�>���p=Y�2 �,�<
4⮈ƕ����x����H�α}
��`�\!�N\����Ē���<�a���p˶ԑ?E�8Ӡ��s�D��q\��8��@�1�d˝_Ê���{��$-��.�.a�>�u�C����縗�n�5\��!^ ��J��?�u��8�k��D!��An���$�dA�)0�acfa��yH���bc����P��_������?i�R��G��e O�o�,���(�1�$wՓl4QLf�Ng��Y��d[��k��t��~��Ö���j|RKssh,��������z�*�X^.�Ur������F}��M���\�i��}�G��� ���ٶ�&���Q1�v�������yZ^�.i9ٺ$�|8S��g8�^]��_ǘ�,Mcq��;��n�o4�i�R�p�VIXy��_�!�ۍ������~ݓxә�5"MJ�(T�=�qcS������֘��4�A�&���f+�>��o��N�x������w����h<��[�®��y��g6��u�G��[~�op��9��>��L��t�Ŀ&Q�h�0mF@��Ko�K��P'������{2މ�����T�>�4�����ǜ5����3������`�px�Gf�q���N��p�d�Z@��P�H��^��u�{�iH�5=�������@�[�PzT��C��^S)�i[&��a�,��ba�i���]���᫓�j6CU���r	�Ch���s�$|3��A��j?���b��MfqO"+[Yf,�M��˨��uV�c����Z�K���}K��#]p�E��Ք�*��he#�o��|I���r�Em�ܛv���C���N�yO��ӀKg�j�r�r�t�W托Y�d�� �.Vfw�����E�
���u�A���Ν`�;���ɒ��@�B�ɍHP8�zg#|5g�N��QPSa��a���T�w�I�Bz��{j#��b�*h��<er%�@��m�g͖���W�{��	���0V�D[\�Cd������
����j 9�:�^0q�JQ1��d�y�C�$�̪Ղ+s�T�;�4�V�z�SD�T��3L+}Q�g�؜�_�M�O(ZT��;X!K�8��hL�f��[_|�B���%��-��D�wp��6m�q�|�j�p�[��hT���$յ�{�����2/���i������ssM��8�Q&�pQ�I�e��4|��&r��#}Y�3��i�� �%�J܁ǜ$@����Q����D~'[MWO	�� ����P�M��h]e����kP���X�eL�n�)��� �'��ڻd͂)�b��f��T��'EK�|g5)�k�[$Y�8àNR*���7��E� :�GexiJ�x�f�3�k<�H�m�Ӟ�5F O�2.�S:Qr��&�I�Ȍ�7R�C�*\�+�+�G��ѯP��L=�!���z�u7K��� r("� 	��dJ�85p-��c�J�x���˫�^�^:/B�Whßl�jKZ�<�V�m�K
�> "�����ԉ
d$FA�� '�t��.����ŀ�mo18�Y�dblZ��>ʑ��~��S��2(}��{�@.������<���O��t�f�wyv~[(��&��Ֆְw��Ct��â�P@��,����g-U�˯+g����&o�ᬆ͵Dv�L��7Ҏ�0��*�GT'����
���L����2�����.cf�8�����Gs�Z�3Ae�b�rJ;	���u�@I����bp��+��n~��*�S*a�?�>��g$f� �σP�Bf�*F�Es��,�E������b���;���	��x�dXP7y� ��j��x���}̠�<M9n��s��y��N��{΀[ޔ77Ƨ��W%��$����(0M���M0���,����H�E����ؓ��|�Wf��|�'���:�h����R�)U��I1��m+ڄx��h�xx.�5nb[�)�Q���i��4�a�+. 'b�@�wR����}�<�%.��s��K�:Ա�ۭ|9�!%,����������F�9>ڈҖ�Kӹ��1�d4�0.��Zt%4���c*��ÒL+;oՌƟ��c�e����Pj��BU�7�=���𒓉��̂�z�(�d�s��p\S#M���O� Ua�{��d�j���7x��俀Z���n��>�]gM�JH�Q�-G-������9�g��$7�E���oi�3������̶��_�(%J�Nk�3�m�δ�R��iT�C���������.�(.Ճz#p���tK�4��P��ћ�3I��D�c	Q��^^`��;iù�+v� ^�4��{f��T' ;�5��[� �ʚ�~�aK,1�*���\��`w�Q.����*D��;��ޅ�������\,�\E�-��AmItH���o�R�;
Z���f*Zwv���Vb����%�b8�^sgכ�>�@f�ϫh�O	rw�NI��!J�2��-���[+����[KP��K�cܹc	Ùҕ�t߸0{B�{�SO*eqߔ�Rrb�>�:%{�iѳ ��[�&�$���G��I��C_�V���򴖹k��p%,nXxҽS��z�?�-xc:*֔��Q��D�1&�dJp?xD�ڶՕu]rSbW$3�.|��P蜨��6p�SǤ�
P�/ـd�b�L��fZ��6+!|���Z�},����>{�C?��E��d� ��V����RG�����*��sȩRUSf����O>Ж_m��i@K�1��xV��蛼z�a�����g��5�<R�CC�v�I��1�>v�!%��k�2[�G���>�o=�w
*�X���F�.@G����#�	�r���S��S*|�h���d�Πn%-�y���m�d�)�_h7W{�},�T�5ȤZ�Q���7c�m��(?����0욭��E����qq���2����N�?�{u&���E7��K}C4A��d���UJ4xx ؑ�ޗ��)�_�_WkO`�vv%��1����%�<6}cq���b)����J�T�Hf�7o`�Q�6����(��#)4T��#}w��Qێi� {���S�����Ȋ`R�#�y˺��KUA�QF�U���32(����"J�+�0��U�ݖI�o0����(�䑀��f��B����h�������t�%X��`R��d�q�Z��N��CӒ�*��G��2{�`õ�V�M"��1	�1��=XnO�ӡh�h B����Q�`v[@hE����w~w0"�&�2�Л.��(�н��my	</��;oՍ�%���Gu����$.C��Z���b�J�l~-��a�'{�`Y�ˬ�Y7��FB�dsN�8y��	Gg$�o��Q��x,GY�e��ߐb��@��L������ƓV2�g��E�>ħ�����Bv|ÅNݏU�O O��G���G��5H=s㛍'ؒ�)�I��5r�2�t���5�	���e>�� v@��OD���`j���_�IXʃ��2ihb{ْL����<�ީ��e�j�����>r�n��Lǅ8[ְT��s��4�p��,
��b�C��uhif���b<ڛ�7�k�`���H1��>d��"����a�a�j�P��������/��Uws7 ˺���qE������N#8�C|��;8��AX⟶�K�m��z�MҶ�{�K�Q��NV���e��^����X���h�I�ef��r=�t��7Ρ~��Jk���N�������Q�1�ow�G��j�?B4s���ˏ�Z�����]k��b��^C��dGIs��U�qF��Cp�ȹ�;���P�J!��d�ͳ����ݏ�ᷲ4Er{oz5X*��+1�dHh�'��U�a� ��#i��."��;�ƹG��͓W��<:�
�Ÿ��ǳ\�y��oiE�Q��QJ��!�
*vU!��&f��q�&|��!6�l��1���6m��B�.��J�9�6��|��U�q�|`�W5�����*�
#��*B���b�x�
[�w�i���)�j��P@��ޑs�M1�.&Vzg�(��͏���ڐ�	{�����6�#�F���%��li�'�ࣰa�,����}��������-��j���>0�#��KqXV�E���Jf~ƹ�
�Y�Ip`�/,��fe5W�1L sZ��1@�0)2���>������#�=�!�&�r[��C�Ԭ(�$��������#}�;=��f�6{S�#WF��'�3*��-�����Yr{�6v��Z�s���tA nd�AW41Z�y�ƣV*ͨ���i�
C�Ρ�lA����CSwi[��o'+����|���~�o�����n�=�n�/�y�v~�����m�Mvl�߭������37�i��讼��;.T�!ʴf��W�S���]�ZU$��_�=��U/�㊕%Wr1 =$�IW�Jɐm C��V�(
jX���&�h��%��Sx[PP@O��h���4:�~�u���LC��G�|;HED�<�/��vJ~�Af�'�Fi�5�b��2�X��ݞ����g�T�k*��V"���~��	fca�H������X�JX�6F�R�1�
�(� ��J��?������X�5����i�P����Rr[��$UbK��]�t�͌�(�m�UdG�����W��7>s��O	���U	��N9�j��
d���g�1#�2�}b��'3�B�O��i�|�V����M��]A%�<�P��t[`1�Z���}���Հ��)Zy�bU�oS��$�և�?��gЦ?���HMʜ��i�&k��Q�ݲ4?��m J�\t���i�}*�bs��Ra��Q��rj�(��A�?�Ck�_���i��[9����v�C}&8h�Z]��MM��G�*�#7��ڣ/}.	f�ꑨ�G	���%� �ඞ�:��;��U���/�)f��ƛv����;����/[D't(��[��? Ċ�,|բ��q�2ޗu�2�'�;d�\~�H:��Vu��1&����|\�~GJߺ�;Uj�g~��x�'��<��RL��?y���̈%хwRF9�n���Ո��Ehޔ<�)�<S����&�f+�ލ��駠3dPy�j?��f(k���8X���L�$����ĻF��d�u�G-m�M�xq��/b��
#M�G�>��yl��$WV��p����e*��;Ay�>��=��I=`7?rE������Z�*�\�[>��kϥ��-��d��8/�c��(�Xe��tXI+к����F�� ؂�(��ӂ���:�W3���8R��!����/��zD��z����9d���j�:t��������ĭ%e��p��z(�*�;koͷd0'�Ux2��Ɵ# c��D��zL�����A��ok>�� ��Q�eZ�)�_���$w���c���N�����Ғ\1>�����72��K�X~�E@�m��C~��D?���^���U�]����I�Ѿ���2B2�������
 ���w���
2�r�1�䱓��0ST� c����Ƀ�9�v
�!H	���s�VTF�[_�t8h�:���o?�qLv���~�j��NM��SQS�t檥���dc����.�m��k���k�â�;%�TWk�dܟXl���_aݎ��v[fFc�����t��`�S[�9�ꑘn�S���jo(æ�<~(��|r����48+엥�˭��$Iu��g#�SH�XV�=h���[�R2;˨?����)⼜'z���L18�K�Z��c�R3���3v8#�4U,��А��(<� ��4#Fbho$-^9=EB鲅	#{���3>��S�q&��'��xN|��7={�,��#�}��. �8��܁hz9m�b�#rQ�ZaV�z,��Me�.l��dK�Qzt�Āj`p�D��ͯG�]�Z�C��~�SQ"��;�ՊQ�K��`�����/����P��	Y�2�\�hR���D ��|���c��d�q�F�N!�qш��7���L��z��Q)�_�{��A+�Dl��+���vc�=�(��;�O!4����뽂�З$U�j�ar-J�`�?r#�T&���_��'20W>00܎��s9Xj(���q��'����a��edxE�YҦGJ��Vu�c����bb�	���������|mu�_�����;���}�b�o��h�f��"��r$���hUuc(��0=oK�6ro�M ܝ���M�1�0����T0=Q�}1o����s��S[�������i�L>q��S�2����-Um�ڇl�=��ct�y�b���v��R\�64|����`��n*��9��H�1y�?z��������W��쩇��g�(�����KU[=S��^1ה㙼A�5����{L\4Y|�򢉌)NMX���ܞ*��~��:���Xs�uL��-�[��w*��q��V7oo��1���[q2���t#cXj���7σ�)�Y3Z��y����dC�7�	������?-5f�p���[~�1A��+ԙ�}�ys�i�؛<@W��箻�G�r�6c8��Ls�X�* �'e��X�pϻ��K���9^� " �!w�ZN1�>�U�M��@����dZ������R�����XY6��}|�-?�����e~?��/����"�j���zN̔�M��rd~:�I�0}�H豔�K{�b��q�c��}�kV��y�;"�j��DLQ��h�FZ-�ͫ}��^b.�+5�;0�6̂ZlA���� �ୁc�il��|�JJ���#��J{'\�N�x=d���k���U��n���mX�]����b1�Zɰ�Dٷi=)F^���,n�!�7�M�ۡRD�ȓ����%�S'���a�Lƕ�hf����Y�5���A���?����X�Hy<o��A�}g�x-�wL�#�>d��l.�?8�Ժ�yO�a�|n�U�Nԇ1W�d�{�l2J�)Zi�%Y6�����?��K�(/�4Z�-O����pnu�l�$�f�޸�-�Ԫ�Y��}y߬���ɇ��2��ڧ�^��=4�֥"��"+QqE�.������A��=��$Ky��JK?\���O�	0O��w\f�d�5��r@\���S{Q_4��rE�#��#��a^�\=p�"<���ak�W�2��o��g�(��pک5��sLn�Xэ��:��X����^��S��p��I��¶Q���{�x1�l�Am�C�p�}������kݑ�4j�[�6z��i�sI�N k�4b�,�p"����SL�3�kO(9<ǞP$\�K	Vs��Q)A ��Im�Q����ie���:~XS�}Q�q�����,�FBoEZ��Ҳ&�/wg]����NQ�K��{L��z�H�*k9�����
��Ov�//9�kC�j{��"�Z�*�1�V1B���<������|y�
n���.>9��I"���	G��Շi��<q����)��2U
��=/�Kz�5[���*����ys��G��M���zǎ�!�����C9�s�Z"+��SlC�ͭ��j���*���������Ґ�g�=h���2��
3i���2e)p��R�bzu�i��-b��Ԍ':,���o?�4��c"����`JM����3�����o��Iŗe�3"8lIr���Ud2B�;����ܧ�+�������v�B��
���Vq?����||�x�JjE��D�F��<�d�����W\bļ����W�}����I-l/:ު3'N;��x�T���1Ϩ��ǜ��"V�:u{��rq�2�kY���9期�O�'�[��P�R�rޙD�*["�ԓ��X �*�������b�)$s����W�������~�
�Y[���ㅫ��^Ҿ�l����0��Q�9�*�Y�	!L����9ܺq�`C�0�D�)�*f2&�ٔ�O�H6ƿm��j��926��j���iR<Iv�������0���[zOG�[R���SARW%ڿ*X���f�o����`�]�8���L�Teؐ]S嬪����
y�R�japG�Wc�-�l�xC�jh��W>@��h�̍�/�!�(w�['g3���1����N� �	�,ѣ��]��	������+C���3��d������h���^C�5:,�\?�p�UbݜD�K(�d�:���N����ᗶ����׭�d�	�We�ߒcE^�3*���ˬh�+��+W͠ڗ��遺�lc��B��D$=�J�lV�گ�qv�w ivLfܐ!�>��\M�s-�֘��| 0u�z]ww��<K����<9�
�V��\�}��ͬx$�Eȯ�=}�xv�'�y�#L���O���k$�f��0��Б:�L�\6nI1�1����5���xc{Z\�W�ЭI���|K[�`��?u@Q[jA�ӑ��.O�Q��'�_D ��o�
�b���H.Ѡ��Ak2��tIDjl�,�\jh�`���,O��b3+kj�|a_��W������.3�g����;=Y��
#�@fzN���#P���{%S�,Z��x�т�_�|��#���t������Fr�-���y��륚Ll�u�K_c��PDG0ܭ�Xe*������W�St�5v� N�ӇB����������S;�H�^
h&�ш�T��v.WO�1�,��>��0z1��A �U��C�/�zLN���� �Z�V�@��ז��~le�����4t�jfF����C����p�=�yٮ�J6�1���c��alݱ�M7o����֝��ݹ߱UJ/L��0�w)l*����d��D�]�o+c���U�����QP�)�I~�t']s�<��*x�6z�J 8����GP�sP-(��BxF�@�o� &~Di�s��1�(��Bf�A�r%h����O8Z��E��M�J��V%�M�ibO&؆���Ga�Me>��,Ӥ&���rd2k�3�O�g��}�Y��l�P�5굾�������Lv��k�TǘmN����i��$�E��QVC��5�'��������+~����[j��DCW����ҒQ��f&Que8��-�Kh�&�*0��E�J�A2%'0;a^'��{��~�&ߟ`{<��S�8�:��bn�{;�s�c��Bp��kp�`r�P�����h�n�ko��]�K���o�%��5妶�gE&\��kq���� _�y���:8k�Ұ3�6��@���qr1*{M�e6V���Tg���u�"�;�M�9t�/�kn.:��Y�W�Ղ>"�5���<�
0�����cڧ2I+���l��38�07`���ç���'x�#*���H�[X�w�Xa��=�G%'�) �4Y�"4_���?�y�}���@7Q>_pN�p�}qz���iBW����Dw�E�E^�|��	�����ѻ����m��1-T\�m.>��q֯-����� ���\O7�b@��!w�|>	[B$����eFH�l���(Bn'��=#�9�r��� ^��M[W�<;_U��[$SJx�1,'q�<F�7(��EՏ�8�Ә���e �M��9e�����,5���Y۠�an
g]1����P�h��&"��e7tP"`Y5tH�<�T���댍<.�5��o�O���ݏ�Ό<��>�9ڳJ��(ޓ����ķ8W �п���6�Z�R`�LZ�����U=F��p4xW�+G�)�I����7k��#[#cA�o�Ã�x�4No�=Du�s�K�_�$�,�b�����G�*���)m{��Vۣߍ����J]sCD�FwCxՌ�q1�{����<��1}�?X^�w�i���q��H�gEF�)c	��\��ݹ�����%��(sH(!� ���M7%h��);�SV��`��Zzs�0�0hP�Xe(�4�`���a���ub��$p�b=������)�!uL��?	���p]ɲ�ǩ0BX��Ϭ�L��:�KH�����RU6�Ia�#�?�~�*�Cn�RG���jL�E��V�<���`��6��Qf�o��d�G^�zb��sԺK�^�4�jl�ɨ�R���Erfe�H����K���pKW����2����1Ĥ�ж���)�Vh��Ʈ'+Gʟ�bG
� �kۄ��^���>r��9'Z-�ϒ��16���)��6@)���[����-e�=h�x!�����Cۚ��~����k��Sr�:`��i5�����Z�RC�[���a�»[���B�RKHb��>��]mK���8���u�!qa�3������s�Sa��X�\wT���KG�?��K�8}�șl�J�A1Ƭ������ #�I�&���F@L�X���"%��l�����TF�5�����kp�h���.C���N�!n�I�m�j3�� ��9/Cc����H����j����l�!-Aq�@�^��ʶt��i���KY����.ŏG*<�~欹(�_���/GN��f����nֿce�-��B�W�i���!� =��ޑ����~W�c����P-!�����"�Q��?�{���Zo�i׉�u��!�}�1=;
t��>)-�5�\��a`E��������*=P & ��l�`r;)Խ� �;_�!��8��vV�?�&���Y�e���r��ZI�����?��[�� =JwZ��D�}`�WR��2��[�-��Z�u;�'����FQ)��L�빓�ji�H6�!?bj�wc��h��G��ڃmݦ�y��5�R�Q�
/��+ii�Mp�d@��-����4���(ݭ^��Ѯ�����tn^�+��Mk�9�_mr�,U�|���D���v��y��-�.��q�A��tTn�E�7�}㙝d�;�Ğw�!J~5���`����(3b�㲭[���d!&���dŕ
���bj����o������˝�1�)єOV�`FY{����J%LB�Z<l0^�;�Ƕ���/?�v~���"�+�m�"	�I ��	�_),'�xq��&�ĳ�6�N����M5�i��9i���kW�( ����'k�IT�t�V9
}�W���Ђ�oZ;�J�;�|o��䬐�Z�qx1k��6e�� �an�C�"+Ǒ2'ǧ�=��-���38�"{ځ�(��Q����^ojv�"j�tS�C8�D?���O8�WWN?�?�o����8�\Y�i�$Q�ԭC��OZ՚��&q� X�/!	���G�����e��7�E��Y�Y!��AӖ53����北�?uPǶ��H�`��.\/z���ώ�)m���0LC�w�ǀ�CV�-@P��Lnn����Nƀ<�P�s�V;��Q�MT6�N�c������R�h���ܰ����F����mJzخ���{��MA�Hǋ�2`Wk*�9g
QV}lGU�4��w��Ki�+��:�������t�I�p
��+ٔ��d]c����χ��c�\7�����u@����iI�~`����~]�u�=4��g����X�Ӂg�9�6/\��
�.���ٛ���p<�``#kfw$\��QG�_5�Pp�u� �H�� �����H�34$x�%WI��`��@�{�pc�IB�x�5/��$&��K��6o��>�b�w������G�&�!�h��K�(Ӊ
��O�5;ٸ7R]F�#�ſp�+.x�s謸�q�ɺɥ�n�Qж��B��>z��={$lߎ��PS���5�%�JD���(d�#@:1e�ue3MBT/Z�a�D���B�t{hR��j ��Ll��X}��]mA�b�f�7c��WX���%mJ�F`�@�f��mP z��n�!f���fW|e��7�(�����K�u�b�\X[Si��|w��_�J�'-�z�c��<
*ʙ��%pEC�,D�2�C�[,��:9���jx-�w3���C�٧�5l��8h��rx�ޭ��2M��䧪��pq��M0�8�����ㅬp����P�)���۞$Fo}_<�Q@%��s��#�S����,��>wJ��[W�F�"�q�d�D��9 �7��f\�
���Ai���MD��ra&(q��]~1��;i+O���a�l�;pq��q�(?q~�ג��x��n܊[����'	A�OJ�+Z�7':6�Z%?i��W�G;���o+�c}������� /�-��t�Ϧ�I�;��ׇ2�#P(���@yR\�<Z���L|Jf��wɜ�0��S�}�W9�|D�'GlJ�E)?����J�o�Ŝ����M��ߝ��(�Jҳ5A����� vw��?*�7d[Æ�U��=v3��H .?���(Lt�����a�����2��){3>����l�4Ĝ��z=���H���)!����ڂ+X���I�؀��rj\��
�N��`Y�6�M��D@��-������	w��]�_	�*_��<0�^{�K�M^������KH�_�K��Y"ή�D���������٬����U@�S90br��7\a*f�Is6L�_���t�f��M�=�ͷ|A)��V߼����_ ,��]"c����e����.�(�Q�@b^��(Y�0����rS�~)��tR;^�t5a:.�}��>��o�Hd>���<N���g �Ϛ��D~r�X�FF�G��ׄ�2c`h����:�x��'�fU�Y�tr��퍖|�XМsy���l���u��Ǭ��l������<�uA������W;g8��?��Bz����7ydc���Pp��J��y��}ݩ�,$u�(�K�Dw�/�'��C����>�����<z9�Oe�����e�6{Lӵ�Zʪ���qs݇��C@"`��\{ޕ�cD�q�6[Ⱦ���ɱ�g�U��9�����|���W I�M��UF��ƚ*��>���@r)�Ş���7p��=[0��I2�u�z�
$LK_שE��:��-�7��������x�{���?,��,��P��[6��m�S8%w{��[܅z`ǔ59�.��0s���;Տ5�Oi���Zw*oa�.Y�Ʒ5�&���t�J�a�����q�B,6��PP�4�G��k�b�}q���Y����=K}�a2��Qk!P���@���j"��\��.}b߽#�L���H~U���;��1�j��b�g�����S'�q��݀��v��wlǄm��gW��m|V�Z�I����2������y�\B��P��E�u����	�%�|�_�̛�R߄X�=�^�ɤd�n>�x�����\�&�BWq�~
�����h1OW�+�f7���G�9���)ŷ��[W��Z}{��o�ɹb���>�˽_�|��k�[_n�[��]UYD��߅L�a.L�Zs{��%��})��S����
D�1f'K^�v|)����z�v	��� 4dE��-���2�y%������}��/e���#��q��תÔcP������N���R��c�(��oJ�% �����scrk�.MV �?���#��N@�7�����$}%5%���H<�Q,?���=�
�u,�f �K�QYգO}��"�k����д�UȪ�����QdG�$� �Bo�֞�T���eԑ�ゐ�(��9�~�;;q�NW�-KW��&��8�/�e�����K���������5>���n���PRz�t��|�[���u��f�q�Ж"3ej,T�#�4&�
<ʨ��;T�H���&V-��ި6U\Hmj}����E�k��^cY����2>���]���ױ�E�P�� �̊I�a _�')G����Yq�j(/����*�C����Hx���q�.i��/��cy][��������į��_�un� �]ߝ��wiSyhё��.�>�MF)�δ�������k��Tt-(�Tc��x+�H���!c�\����V����:��4�kg���1��o�Z7����B�c�QE��1�%�SdS2�X�iU^T޺�����M�e`����(���J�}��ɓ���V�0Y�;�Ifv��+����y��:,�{abr���fCM�&~i���9ԓy����Ν��kY����:чZK��χR��v��x��8��Q>�l�#���s���I�`��IsB(�vR���D�OglT�V%���x��{\t}5f�*)�L²O�b	#$N ,��k�-��;u�������]��1ԝ�H���H��N��UI�q	��6[�u��$ѵK��8�[Eyh[B _ӎ�J�JC=m��C�����{="$�B�"ި�v���{G���M ��	W��;qc��s#��A��]D��*L*¨��k�n����۲Z"h�%���΄I�i%e�W:�s�3����FSHS�u�����c�� �q���F���"��d��MKl����t�EM`�C��L�%�b������sU.
W�>sj��+��p�Yit���	�
��Q��pkm���N#�&ic4�ĝ�z��Zp�M(bʨ�,�V���@�B��m�,]+H8ȆҒ�qvHsY3�.�,=�gup=r�".%Ib�ȃ� c�xj
r�G��N�s��b�nZ�# Ŀ:�.J�K���|�迬4��#���ST��ҫ
ь�Fӄ�4��/_�G��΅S*���HgSF?�;~'0e؂&#���	q�8�Gg.C&~F(oW܃a������A<�|-�*�z��-�(�0t�%t���;��A|�������Rݡ/X���a��2����fn�}�������g.�,������P8d�f�� }9Wʏ���t��ų�yZcla)�f���h�������O���V��_R��D?s ���82f����x�x���H���jҟ� 1���N�s(V�?@s�~<��+��N���
�NqQ�R�$h�ƛ�9\kD@��-/9��K�d�l8F����ǅI��E�9�"��d�)�F��r��.g�pJ��C��b�%m$��;B�ډ�)W��
�#�8g�
%U�~R�8�*|���F;�HГ�"��fs�}U@QG�U��á�v8�5�(/*�[�h1݊cQ�P��8���D��]cRF��ڵ�Q�8��`A�Ҽ-ǉ��~���,qlͩ��-*=���2���8�7�׼�)�_��������=��-3"�u��(��|[��gҬ�)o��W;gk 08�j�)���cT�o�t�F�ΰ+b�*޴.gu��q$�B���!�$MJ��U i���"�w@��<��.>���	�N�.���x�5쿋FH�Yz��#|.Eai�b��Lf[�I:S��"]"����5m����'�=6��A�0I�7�J�	��؉$l5<=����D��<za06(��g�tƻy�f��P�a�k�d#������S�?�0��L �x9�%<����&Rbfћ傮

�~!ł
��;�K��Q�tly�We:���haR�'3j���5�3ioϞ��4�W��,�n�Xli�fа���G�>6Add�$���џQZ���ρ#|^��Ct�ĩǿ4P�@v���F(f������S�f9��Ҡ���1��^�υ�&	��<r�8�#���J�g�f��RP��S}�����}k�-��f�K���Qb^�6dUi��f3��(�gg*����!�����i)�^��g�Ԭ.9�Z�[ߌ�Ui�u4,%:���G�Cˏv�Q�́X_7As�I�R���;P3^��({J:ii�_���>�ἯFd��k�M�ͥ}��N�}��n�qE�'��U�)`+h'i�d�~��f�,~��
D�G{��Gu>@�>AB�1[�gY�s8O�ն����?�n���;�_%mvc�-'J�D!X�v��S³/��j!b��O彜��!�Uh�p�?���,9���E�`glrbu��u�ٞ�1x-S��3�i$�g���dH8���P�}��so� �ֱ|��?U�����R@`^?�Vo2A��i�mBl퀮���o<x������;��R)��j�,���/�ֹp(~��y�������LP� DN�!璒o$�.����O|b��[�mt�[#h�ky�s����p��
��L}6Z�%Q�}.%FɋXg�ɤ���k�qd� �8�_���	����P�u�?��5`�Љ�+�PD�83�/	�U�����f��7!�+��a�ǌ����n��Q�1�?y��80uvy�)NJ2ϐ�r�Bh���S���o��s��} ���nG��]BF����{m��B�C�A�ծ��u�2\�W�C�f��|���%	��o�e_0���>}�%*z��M�Z�k8^p���=-�np4�F�UDԒB����#�Ѫ���r��M��V	��o��Z:�dCn�P��̠��	�Fz�� d��fz�Q�O����t�;T�^�%���D�бK-a.%�ԑ�Qaa� ���̰Ţ���z�qH1��,���Np&���`���uT�c��'߫z#�v�lo�l@�E�C%i +m  Ut���/ޓ8�h��વ��E�96�N���� \����9h�őp�m�G�BZ�g�Р�@���x��Sժ$�x��[�f-q٣0V�י	#I[��u��J���cA�$tyvbٴP��U��mc>�(��c��|�u'J���)o�k��?)>��=?���1�-vy曇�I��'��,�}+V����:w�-�wX#��Rz�m��dvq�n3��N�]���*�22�o6��Q$1�M�G�1.:�)�/ۿN93/���%z)�����.��L�-פ�K�W����*�U	$�c����9�� "C/�G湀;�b��)8�2װҮ�Z�1�߮B���n=��Ê�x��O����
;��q\t8����PX������ZjJ��J���jº��O.�H�/��f�b�j�	��c��T��,R��Rn�����8�7R;f4%̡H����K������Ә���B��5X��u�� !��"I���*=�D[-��u7�Qc�N;�����ɍ�d�V��f�
D��m���8�W1�]m,�	�"h��h1�M��u(T&N��fgH�|���-��f���<�
�l����]��q�u>gJ�^@��ߩ�C�[�7�������@X_p6�U �~�kb�J<ZF�i3@6!���⿿� )�;�'
t�+�Z.����χ*3^�1�����.f�m�<�t�k�EWr����YѨ|V?���{�^�X�2�^]��
BT�e� ��m����Χ��C��	�ƐT��	<�$=��� q�l��91�-�X�%P5>P���r+�Ӓƀ�^T(�'�\f�ߣ�Z����	y=^�G���ؿ Xq������(�Ex!��S�d�7`/۞�l�;�� �?��6�*�S�Xx����g�~#AR+d�Bc���=.%�����]�VD_8k�����Eoa�Luj��=�e��������bg���{kzn_�݋�-�����f�q]�V�"�Ft-�؏�gAq�X,�r�����^�^��UN��},9��<�z��3���_�8��BC�wEnܑ�.d��<pΐ$9�=^�n2R~�<���E�aN+�p�\qE������)�I��"G��V��S2���^�S*E�`��O5�� 
(�=N"��F'�pQ�:�DO=��a���xÖi�a�mE%H7k]��sFG��n�4��=�j�I��N�
1�N�Y8τ/0�;T5z���2xE�q2�	�V t��P�D�eès�FTY�� p��MI1%F-^]�8j�������ε�����!׃�I����e�����=��,�I�*���4o�K�����Gci�<�:�����3��?���Dj`
,X5}`!���k*�%����U�ܸH`UM��U�u��oC�}�l��o�ޱ��G_3	��b��G�2\/�Q���f�U�f��Zu�r4� �e���)C����{9���^*�C�+����Ԍ���o���c�*��݅��T+���݊��U��m��j�c����j��ғ�ߋ`�h�ICdݩ�]m�;ɋͱ�Wtɂ��rk������2 d�U��z� �� ���՝��Ƒ��aMDk����jU�b5sj!���-f�q2��uLc�5b2���6��M���5���a���:S5=|�Ԃ��8Eĩ�\�a����9�x�W�~��閤H�����Au3�԰��D�`O�{}M f�����f%��Fo�۩��µ��M����4$�D"��2M��MOu����y�QcUN�^_s����������%�[x��̈́�<�Wh�����)t&�����vqd���ж/ e�^�h
.6�� �P
�[𩷩�M���M��K����9a(4u�R�[��0�9�뼟�[��5`e��[	��QE�E7������j�	o��V�>�]_�JW�����=�rc� ׷���80�`���!�F���!߳��n�0qA��t�f�xh
a Ԯ�j�`�ƹ_-t����8:
�sD�g�'�iU}P�'Rh���<�ު]AN*;0��qI�5����͘5_�x���<)X�+6�E�J�k��\�A��Ǥh.j����MG~��f��f�?�_�k�\���:��?�O;P�^_�&ѡF��ؕ�Pǖ�g`eX�����vN�(J��� _ǜ�o�Z��.l���J����õm��܏���)���$Lf*��UZOZ�6�1p�͙U�L3X�ڔ�@�l�j�<�7Aw̿��*�eI�5��F�FK�Ő����gTX�K������C_{�|�9���Qz>�� �Vh8�;��gf}�)6��H�����x���6ֈQ��Eʄ_�u��7�L8W[4�9��h�a�Zo�o݂ �h�����&C�hmd�+d�-����}����4��i�q�)a��A2LB*�V���cKC��z�,ki��qL}�k%�js�&�D�{(i��Յ*�B򨿟�.��\S=]�u�{7���9�'�SK���q��G��vH�Уw��`FJb##Jl%��IVYK)B����z��m{�O���ImWHf�嫇�}����ݮ��CX�,���	���v�
���8H�*o�z}>z ���1�*�hP���}�����l�z�l=�L�����%W���a��0� v�K;�/���@�Qw�
~��\��1
r������͊� ��h����0���k����.��d0�Z�c�J�>��Sa/��k8_3������Y����V����6c!3��Xh��['p�!p��/l]�,��5��D��_����&Iٜ	�}�L�仟���y��1r0�1�~>�\������Kete���A(x���N৤��0�������z��n�&)��ez�t�W����e�>?l�G.�V�bD�'�R�aҔ�v��
��Cm_h����2A7��V��:�6�K��a��>?)&�,l�Վ�B
������j#�֋���aS �pU�%�4ar�ieR�^$���m>ّm���͆�v�����ݔ���3�n5j��RF?��*�֞ңS<��}�t�AfGD����sn@u4n�r�o�w���G+9B|-�y�t����:k=��Ȑ�~}m��R);�&½_�[���S�2�,�by��E�Z� �Z�1�����eO�O}�'	��^�M�(f��}�d�4�b-b#��+��ȶ�t_�F�T�'���Pt�N�-2$�^$�Ȉ�IL\y����'�=hq�<�R��}ge���sTVm�HPD_�ܫL)�z��ˌ����iE����C9�\|� E2���P�!v��I�!������N.j�"7�W8z2�;��3��r�m��]Ƣ��ʚh6��p��]�"L��C�j��ƅ��b��d��$~0�����ﱫ��+�����Q�\юd�_F�m�k�U�fX딌����	z�{�8���]f�z�82���|�A{E04��i-�ބ�jp�j-�2�&&z��|�G�	z�2��~�>��\��@v�aQFr��dr5��H���f�*z.�me���(tOC���:�}!3�&&i�����H;�OU~J-���o1�S�G�H�;nEU̫�0m�=栾�P+S��um؛�n�%;m1��4������'�@g4sT������C��f��Yk�,��ԏ�L;/F;����)�[�g�J��NCo"���J�XW%k�r�s����E'T܃�������yov��̞��f9�Tk�t����[ |jm���@>�U��6>Xż�ϯJe���i�U]������K\7�Á��uC��t���;�.ww��c�+z �X��a总�p���R�=�R$>��QL�B�uY�������8�G�����|V L&�Bf�hrp%���P��\�b����BE�y��nڹ��4��D���O�Z��`��?�m���~)1T�/���?nL��( DD���el�0^l���#� %��MdJ�A����>�e:w�F��ϼD�ǂ�׺����KJ�㭘�y��0I,rǞǙ�`���Kd�blO���
Z���FgD����~E�,�
�$"I�p�S1��qq4{�3%���+=I ����N�*濝�YAFTf�G�#�%���g�12���'rN�@��#���N�x��Z&(�Jf^
q��C�#j��Y:"�z�+|t���Ϳ�����xH�Dߓ�U�N�j	��XI���od@����a?�vY�j�I�Eл|A��ͫ��?9������]����8x��~����ΐ�H2$а\{�Z�X}��1�ENI���-o�!�ǆI�)���"��J��=�<�G�*���Q��4�B.�r�/D��O�~�z8�f·�%%��JL��Zz��5ټ�5Ϟ�I;$.=V_�����hW�P���p�+0�.r"�X�ԥ� ������
,? �h�k|����r�&q�(�z��s���C������p	R�\�޸{�����ut|2S�𲉝�����Τ�^Ga�;�����%����eM�U�g*^�J� zӈ�$�xY�֑v��*�������c���*J+ٞ�A�W$�z��+�U����WJ�1�7��	,����:�\�Ջ�gyh;@9�%{_������nL�b���h��ԞB>�����v��B�]7_�܀=@�Ѵ[~���vں�~Z��IC�E��HDL��%�(h��4w}ᷭ?��~� 4;!�	}L�|�PW�����z�� �4���[�{%7���E�H�(�*z1�`�zDn�+��G�CP#Z�x}��z���<58.:Խ�dY�S�E��Bd�:�C���ʛ��E�͇�)�|�Q�ĝ�0��j�S\������x� $�zy��
 ��Q��U��{�����=8���|�`����&�#�'H7�갣�WJ�!}$h��E%U#��0��b=�j��ߩ��^?�n>�9�. \2�e70q(O"��ȵ?�s��3&��s�iU�=��i-~ځtKk�������
[u6�Ơ<d���\��r�j�ۏ��dvUVޫ�Vhs#�(��U��}hL2���v/B�֟����@����<;R�:X%���f^}�C��3���&Ws���"�/<�1��`�o��P9� �w#���
�-V���-ŉ��E��טb
�w��FQ�Ь��&�&b.r6�9$�Z��m�����?����A{l0���*���]�+H,a6��S��n����v����">�L�fƁ�;M�!�@�[F�<2Q��+�����O�_*���;���v��f��K��t(/�f=3a���� ��j\�)�����K�Ɉ��F����_�Ӌ�1�'uy1(��$5<1����mj�G�1�ĵ���+���_̿��{0PT;���d�,������3��.0�o2K��tc~�m����Y���s��k��ǫ�n��+���C�\GdP�3����$(hɅ�x��~(j-<���^��;wt`HtT|	~�,���6q�¯Q�v���z��i��-����n�Rm>�[���V��K��.$��,��$���;��E�U:��?p�l��֚������}������E9���JsA�#"� ���`7�X�+��%��L*H��^"�v�{�0M:T�<�sԝ�h�Y^����== B�R'h��W!�Y�(��&j'Ţ�W�>T�5v̀@/dw�+�6"��Gh�����2X����c��ky\h�u ��M}��0�TF��|$�� ��[T7��� ?�6�6w�|b��½��	�A�//H��M�,��6�p���}�hr�]�q�9��'z�e�p���>pZ;���ѩ�d�$����̛�.��3� �m�N,�&,�����_9l]Peu߂B��?�c��H檰<�B3�/��6�����mt���s|"�^�нa�P����sT� �j���x���� ��v� �=p,�IZ��3"?~�Gzz�J@@<U�\�bs
\[v禍�����x2���HY��l~�V}�X9��4��g�
hi���4<�ر�fY�@9�*��a�QAi���j�y�`,�/`o�ڵ�N�^4��z��WL �;-0r�㭉X���V"A��b�3�	��H\�HV��_#+�ґ[U@�#�����wq��|9^K��9�����w|���ٗ4��ޚ������zR.	���g�0���(~�!R���|�9L/�O�b�?��oa�ywfE�X^	&�_��qH�dC:���Gإ�n��DF�u� �����(��Q R�.p�ƸD����3;���]_�n���5��F�+xC�x�P������G8?o�۰�\�`?�WMo��ow�SA��n��<dM/�գ�؝-�
7���	��Y�I��G����+Jᒁ}C� �D
����`��I�I�]�q��Rf5hXKK�$��y7}�����Kl��7!Lf�^mG�r�|���?�hwW+ҥDKh��@�����A����e)�y��)�/��1��-%����:�^����;Bi�_���6HU����èC��Y�埇#���r�� =�%|S�ʪ�s�;����A��%����q��`�p�?u�+���l	��}��z0H��^R�X^)�sKhl����	{�P=�@���9���|�٦,݂݇��$�Qm�Oߥ�`�Q\���5/�D�E%�8��S%�]��\q&�;�D�|�

w�������S<��ҠyeAFy�&`@�S����:%�yR@\�������׊ֳ�?)*Ne�F�ba�e� b~-���:k�q�$,&f��֛���%��y������2=���٫���_����r����T��	�r�c�c�)V�f.t��b�١K�7�q{w��ق�Z�PFb�H�,�B �+�k������s
f�*z{9P��-��%1A��5W5��;�ma��Ő%sz��Y� �o����z5�	]�UR(O)*.휃P��nu�֝�ک:���L^n()f�e9�H�o�m�����b�^�`6��8��P��F�Z��B8Ⱦ���O󤅖�F��8�_�l�W��&��yh��?����k K�/I�"�#��u���u�����z�Zt��Z/'���b��y��2�\��7_�EfM�'SY��ܺ����.�I"�{��v�]��"dw���l��_{���K�}�� j����y�DL�*&x����DnI�x��c�v)�F�GWu�����jڇ��jD������@�`u>�^�c�Ao�O0��r`²^#p�[<4�T��{���|���q���B��L�k ([�hki �d$j���`v4��n�Sҵ#H>��ϕ��j}�h��^����C�8z�����h��L6��(���Arn#�k�b�8m��c��e؏9���I��������N^�DVѾĝ_���7 	p�(�w #�E��^G�#����� h^<W�J�ջ��@��y�H�Ge�&2����Qn�7�k�g�THŎ�C_�8Ɛ`����7�b��[7"�=k;�^�>��/o�V��ۅ�ᬰD^HSp7��ϘU�>��"l��0�p1J��RB	[l��1���nɹ)j�}�,;n�Q;P�+< ��/����es��U��g�Yk���xk��g��þ�2�:gQZ�l���H2Ţ�ެ��l� iҹe����1��zDB���F
9�'��/�
y-�-юVz_aj!����� ��
���׳�ˣ�I754��aG��Y!S��D7�<�����C����&�%+�$&\��y����U�1.��5-�*b>10�TsB#�ͳ1�1|���_Ɩ#éǹ/юy�K��}^��
��u��j򽫅��(��y����[�9�pS�B,���hr ���!���;����k�Y,��"/�f��r/	�V0yu_�'g��KH5%~Y� ���^]t��C�F��X�|X���Q�-�뮇:�h����P��r��[ty��=�^i����%�I?�
�w�(��s��K[�p�K.�O3�yj���y��|��g�Jm>�x}ѳܧ'�q��g�5"#�{�k�L��$+Q΢��s��6�8�oK~���������j���j`��YP�Q^E���*0+�m표rE�
�4,����.�/*����RK=�k(>�nr��lw��-���p�6͇#�Κ5t�&��	p�K-0�VM�f�P.��:�b�	��=��^����{l����gV��|�W�OgA�q�K���0t'Y��C�1��(�a�N�q��s�U}�s���s�W��˴����Ϧ�k��(����UG�J�kU��q]����Y�%BH	�c'Ў�<*��/C��-�h@X�).�1�ay�3�c}�hW���òi�z�]��T��"s��!���~'�ALߞ��|�ͫ%��a�~�(�w`=������֏����Vh�܇��Su�Z`�NZ�77���������v#5�FX�!%*�+��>��,�
#��4���Ӈ��UF�#"g��O�l,�!6�%3���ځܽ�@&a��0%�����*�z�}�c�#첌x9���Y�䑕���-�����P��y?�F	2;�j&�-��;��%Ƅ����Y��1�菜6'ŉF������j���h��#�X�m���@B��������1^�+P$�OTo	���z}˩b��D���8�����&�'^Q��<��F&�&o*��wt��P%�;́�J��dc�̕�/)ߒ���V�&�`�ǆJ���[�� �/SA�xc����7,u�F#�JX���z?(�)�4
����������9]��1!��A}?t��oU��T�v8���1�[,�/v]�]�X�u���_��/f}㞢�^ʘTR6�j�{D!��v�.�G�M)��`��U�:�������YX�OI�>��'�yh���{��Q<�[�'/��n�?���	�!L��5뺹Ñp@��)�����`n��Yud�u������*��n�����FP��;��9��B"l��_b�Y�8��S�ݞ��zC|3G�[�eo�J3�7[���Vr�X�s�"�Z���:�SSL%������y���d�J�R��Y>6�FV��p

y��4ޤI{�M��;|Y�W�~�J�D��WEom��K� ΕJ�J�yǧ,��`H�--�^�0{2*u��[	ڌ��}�|�C�����z�M��C�\����A�Ġ������ʺ�!����yhm�G��a�!�
��-r~l>�`�A��G˶B��� �/wr���`����N�*	�Ǵ�Ҧ��x�=Ԅ$[�)�&�@�_�"������D%��/gGU�Ow9�>��qi�l�2/��H��EKNx�G[�yRK_���b�p�a1�?3j!�0��2�f�(�\p��r��ڙ��7'"�C�-��Ss�^]Bx�9��I��F��������s*�%�׳jVĸg4�jL
Df��^�?�Ng�٬���� B���0��KVm�����:M:�y�Ko���i�]��D��-!Ӽ>(��׭�\�M� �@|��-ߨo�J�ګ��=U�։b2R����@����,�*��8�Ms&�ʰJA4W�UO�����%���3�r�\��J(�F��XJ^w�$��m1�e��b��~N��x��/W��,m�)^�S n<O���>�g�8�GQńI�d�\z����Yn�5
�(cM˫�E�����eR2���id��/��u���A<��l�tWs��~�A����$��@�]�(ʜ�/��{����[Ȣ�o6(���AB}Z��[�|~rq��f�����-eI�R�����m�ZѴ` ��;�2�_B��Aq��/� D A?���#���e���Z�UFNȴtz��6���[���
�il��aأ=��`66���7�5�6�E2���[:p�1���)~I`_�1f�Lˀp>G�`�rQL������X�/~���L�ZΞ˲�Ũ��i ��Z�*�,D�~�Õ�g�)����^�3a�E����6$�&��g����w��t�W�xn=�E��X=�*���j�t§�y0u�u+�'l�Xi|�? 0'���c�����\G��y̶��r��շxV~N&�1���塝,�w�T�>�^�B͵��$�z�fW�$λ�1�>)��<�O=��bWBC��j?���s����.�yś/�W?F�ְ�\�0$1��'��$����"��v������sQ���%�#��B�MA�ދʄ�pS��f�Ï˴C� F ��	:=���݊�d���-8�-�lg�sW	j�ГEX���w�U�3{�����9!�`� g�C�(��"b���eU���C�+vw&�<��c�P����玾>g�{��Jܡ�ᡠS�g��vU�Iy�!|���P�����~ �����Z�Y-��� / �,��2F��̙�kaA��V(D���j�qGym���βu�JDs�k��-z.:�2tEU.m ���i\��Wgzj�]�����cͅ[�R-��G�,�Z�%Ѐ�٬�7�Y�a�,�[�����a�v��;�P�ՠ-4������;�d��̊� ˡr��>���Zg���J���M��G.|�y�� ��֊�ᚦr�(8u�(���}��qv��X���x� (S��so:�R�TnDT�N�+?x-�
iD;;8���$R��B��x��H
�f��D:ϛ*?tN��uop��T*<LH�����A�PVݟK}�C�s�y�-B��c�σq3M���8��|��~%���g����>��	p���Q<����tӾ�����V��`��m���u-CVY��]�Wp��V_����%�$%0v���H暄Q� ��ج%��n���J�r�&s��R��}�`�^�j��B6�x���]�J�R"��z�n�Y�����WK)�	m^/���:�S���`� �Bİ�tè�R�Q�6��g��Y)R$���84� �]�x5��%I	�`�Z;#o�;.��;֢66�?����զ���ȷ9ҳT%5�V������5��*�ݪ�9��1�$�!Щk�P�_�u]�l�E�#���$��������8(D[nT���8�J'u�܎�#3���0qwT-l������7����	asAt�|�d�EV��D�9��]��O�o�+�u��'WG�^��^���K"���@5�O�����Ģ�����]arH�Ai�Z�'�����WM�π��-��>�myv�1��q��
������o���m�������	 ��ۖ����&;� :
h�����PZ���U�	���^@[5�Zs�C�b�l/j��!�J��6n��ƘK���'��o!����:-�x��(��Oe�*�I}\J �>���,!#m���f$	S2���HB��b�WR�c�lB�z^2v�H���gL�9��S��-_����D�z3�T�-@z�[����ੇ[[R#I_���j
�m�ܫ=ʡ�MSyi����͑���S t�vId!w����	3�a�a|r���X�v�z -���;�+n�����qڸ/��x�)��F��.9؁o�����H�)�G#Ng;X��.�B��r�x�ͼ��W�Cs�O5�kV��:���cv��d�������;kVogV�Ew���І�{;y�TVb�w������}�S�?�Bԉ���^c-r��qu�������rM���8�n�,��c���R6G���!gC�� "��x:��7��t¾6���/DJ}e��M��MZ����e�9����-"lm��x�Q��Z:OD6��4m[�|�wH�i���}$W��_B���g���J��R����� ��gN�4��[�_n&���6I�f���1kNG�H8H� �}(H�[,�y��5U�S���Nx��Ɇ�n��l,I���؇�lz2	����Þ'S3Z$Uk��Ȟw�d�_$f�_���.������x`�Y��y);��_�g�FX�����x������x�f�>U59�ot�xl<Ëyw�hRsF�do|�#�'�=��S�%��3�YP�:Ɩ6�f�y^i�u�H���X���R��zR�b������Ic�\��O4�I7c,6���ﳠ��H���o�P�U�C�BG4iC3������-x�)Ϟ5���5��,��>&���]�3�F��U��&�R��]z��ޟ��R�Y#����W
2C@_5�(	��ӟ8/d��՟��>�I�t��� �?�����[�6lC���q$<�'�߾EV�g�"�F&���~O=@�]S ��I0��P��/V��Q��ⶤ���B��&�g���Y�X�0�@�B�_�m} �o���*ۇ��Ne�׭�F�w,�ڗ)�Rj�ZQ�g�GC(}g9�j*�g@��S;�Łap�f�o7�ђ���/p�w���F |��H��y�]ϗ�z�\��;䔢�ew1N���

�! �
�/�#�4{�E{o�eG5dp�A� ��U0yiE��k���Fo$�1Q��S�^Mb_��'\Z�����찘�����(���3�a�	0/��zPʲ��`�c�̌TBD��έ�v��Q�a��&~j�le�`)��y)pY�F]D<bCb�@FC� #z7S��h���@��<���1D�h�BC��N���2���sάln���U����:PJ�ڻ�K�&YCc��G�eZ lD�����lk�������ų~2ʤ�3z���6�y;�]�t�T�- ���B��Gօ�Qɚy�� ��������T�~��Yϕ'�`���z@ġj�+~{��2O�nK�e�5!� �����2�6��Tߔ�͙#Oْ��� �|��9�������o��J�FD����Pg��nj�i��[�^ �௏;����@8[>�D2���=��{6]�����m��̈%8@ʩJ�A塾�*�(+�AI�'m��5�Xk�_Gt��R�s�%je�me�g�\�A�Q.k�'���}���!` �<��4�o�O[Hh&i/�%O����2�dwތr�O��3�4S`��+��K���g�1x�J� ��_�K���m���3A8֟
�����|]T%��%�mD=`i��Dƀ�[��ˊ�^sۅ��a�X��,���������Pa�G��^̥�P�@���ӬX�����p?�*����cR���ܢ��g�ōS�am�Wzo�;4�ڈ닒��1�Y�w���Ԍw�}�$O���ϫ�y�����T�B�t
��]4��+a�}s�-�����*��q4E��]�'̇*���1L���91=a���ч��� b~��"H��b��mt���d�x��;�C�&��� �
��p��5钿�0y��D(b�ܹ$P̬1��%���)*�=t<3��N�����rY�WS��Eߙ��@]�Y�5U7Զ�p;Z��>�=����6�s�5
���Bywd�,T����a���"��r��K�SJ[0�J�%p��/�{$��~�[�SiU�j{q�!� $�rKV� G��E��C$_T�8Η8�}�5���f��$v��}ɥ��[B��|&.m4�VV��T��Ô���Y2)j�Pi:@z��M�d�~��<Ү��?"�2D��O�@	��x�س#OlBw��vB!�ꗟ�%�� �7���N��ñ��<_ux�L?2C�p�r:��9��d��Z�<v���^&G�j��3�#+4?K���F�ͫ�~�쩱P�C������*z�΃~�$��4r$��y��]�;,��1ů�~�dַ�tZ�?_�o)ڎ yF�,D��4S����%�X���ah���,�.�;[�GPG�ǧ�	�,�:��T����qmZ/r�}$1-��~o2�:�*����ؑ�'z=,��T��{B�����s;�t]����ֻ⡽Ί7��j���((�k��1��)����R����͍J�_�Nyu&"v�X-HI��������J���\��]WG�z(rJ�N(��m=V�O�^K�¶$O[��ܹ3�j��iO�d�@����GO�,o��B�#X' +ŔV�*��غ�=��?=��R��[ab@x�s��M�ف���o���c°�P�+svq6��8 -�\[���Ϫ�J���w,~�ח��	K��+��*���{�����3�v/������Ǣ�N�����*à�z�'��8Z��o�;�V��?)�Y�=�0.��x�w?��W3�ۇ������K|r9b�zU<;z�6�b�Ӊߚ�o��zs�V]+�l��XD�&~���n�P�}yP���3��<)`K����׊2�����Q��.��sQĽDO����e86�Q/ ���˒�ƍ�:�[�E኱�K_�h�j�bm�ˇ���ӏ��w�)�\Ɇ\���pg&�"���?p���8.��-F�B��p��H^�gⷀqΏS3jaH!a�\!`M����b��qu��h�`H~�X�����u��af3�I�^ С����cJp�E{�;#<�١����������y�ө��b}�|%�#�/���\D¦�!� (�m�R)�F��1�(����@Un��]���o�gJ|�ވ6�S�W�e�W�T*5��*���{]�c�ᑖ����ܝ�-�O'��C��k�A-A�'!�]F�l��%���$�=mAN��[����� O�U�٫Bφa,���=�n���?O�8���ε�+!q�'J:G�;Y�tZ`!E���2N�Cб��)T���k���ޫ5c��KY�����w�9}a�����&�!�n������/+���:�^��Qz?���]�ɍ+^f��=�den�ȯMq8���+\mqbk`�-��9��M?�G�Qk�T�TR���")�袽���ƌtF�c#���T�8�I��>>�c����d2H��i���-l\��B������4����;E����	)��-	�Y�`B�<����)���^ 	����U�����%���<2U�{��/�^Ƚ�.f�c-H�F��H���	P~�6:t�?L�����{�U����9��Q��0���c��������P�(.3m�����H�]G����DӨ�
��d�mE Ǯ�xݲ��(���"�!��Aa��CQjý�G�lo�G��N�9�VU���/��+�o9	�
Db.�e�N%�֩2t�Ħ�!'J�?F��@�v��6{��d�ڤ�"��s���h��cp��r�S�Gz��~�@�R�� �q��	��6�w��R���J�	(n�ro�.��=̀ۻtƑ������?�҄�k��L�� v�'�Oj³s���x�>�5��7�#H.�<��~ymS��F!)�gIʁ�F��hq/�-U��eτ⼍祠�J��"�*#�2[��=͹l���Ύ-$A����-!x"	�c��_���k	a%�s��Ϝ���8����H���Y�chh�� w�q��C��&ࡥLբ� ��Kdl+�?=-߇�A��+��=!A�����ݟ�	���:ϫ?�BuR\�܇�^��8�L'�#`3W��-L�Q���3IG�������#�5�w��W�}���$��.���3�Ί�\�}vr�^g���D#�L��8�Ѡ�a��7�|]yG��2|q3ϛ�i�l�#�K�$��q0� k�ڙ�ؘ��P��F�5�_�-و�C�[RJG��a@h�S���'1�C�ut�L���)C�lhn���#�^��ȓ�c9�V��@8�%a0B ��A@���<dQ<����<�^buW�2.��[�VL��"�&��<Z9ƊC���wS<�M8D,Ǹ訣��Qh C+���P*���8����y;�2}� u��1`Q߅G��+�����ǝ���&j�^�/y=_#�	��:��O�y���f����c���ݨ��A2Dx�0�!2a�F���^f�!���������^��dS��Pl�
�
gE��$�kf�c�2Aظ�w&tnn��p��`�'��p3���p �/*�yB=_�#�f��s���K����'��'��iO��⏛}o]��m 8��%�A�~84�)���s��,�2��ػY�lǽ9��g��0��A�����q�1u�v�Dy	߃L�d��6�:h��,�mj�0Uʽ�Ƹ�����¸��<���_���n9y/�n�0�M�{������� uՀrv&g c(�S�LaR��5�㛻禎W��7ӊ��H��������PD�8�;S�����g�H�xm{���yx��'b�'.��r�P���3���&%��C��t_�{��'�.���JT��*���W�O*����'h*t��c��mc��D��o"��Nn��Z�;[m���Ԋ'�p$�Z���t{����i���1Ds5ww�@�ʽ��麜�t4�D�U���*��h �����X^@�+���.1��k�<�_k@�.��sm�)�H�w]C�8k�Z�o�s�G��J��$쿅�Y���0S:�����AYu6����h��{6u�!�sy=R(�a��x�\�4�ȇb|��ھ� �Cg�%�K��T���%���C2�J,���r�H���pn�s�q����3�ZG^�e�.M��NKH�$��S⌮���pJa�g���]�,HTW�~[Fգ��0�r�V�}r�i�`��+�n�#��9W�����HL�RC�V?�����[�2�r����A�![�����,@�)����B@�R�U"�C����f��=��z/Xe� &�6
���	j)Bp���摸V;
��<�4����f�l%}�\���Eb����'_ĭ�jځ{]�|����y�W*�ڏ�j�/�7��O+�G4is]��9���)X�*m��g&I������z3J]�4� W�^"ի��{y����?~a7�ً��Ko,Z�з��z�@ɵh�6����PYe�ͩ�B�#9S;&�`���$���F���E*�)��
I���t��9������yf!�] �a՚@�B��l��E1�����a N2�;��Hp�>�������l+�?�ȿ���=gȚ紹b�����:��L䌇���TO�zׂV&�,�����ӷV��u��xgc����w�k�(ݶ���r�+_g���x���߇[�)oޜ�7)H3���ae�?�s3t�����lOUDF�3N )á���TqkS�����8oɆ�����Qa����6�#�A�d����q�%J(�滬�Gg&�5��1��ví@!��{��8jp�D�#}��@�qM�P�~�T�(F��cRV�g�o��Z���H������W/jL1��{�J00j��J;�ԭ}��P���w?�����5[~oKX��g�� �����pRo[��	�j_N�8�kb@Rue�*D����w/�eM��L�d�8륧��:c1R��`x!9�b]y=�o�@U��&�V�0��T���.��2NK�k�Gvy�׆���ӎ�[v��_"�ۚ]
�-�Z�(�eV�A����@����R )��NA{)55����s�R�W�2I�w�����H�L�'�� �|��A�]�y���[�}A
|2��c�n㗣%f�k�=���.T��;Sz��#��B�4�zC�ٜ�?����A
�* ^ݚ��ݙ-��ѧd�C�� �>�q�n�>�@b���BW�;�Y"d��O��Ɉ��d���w�x�4y����
�	�'��!�Gvj��o"�"vG��v_���k�m:
K��)�2�
o�M���.8�z٬�WH6Mf[Ȧ��J�d�	T�I�ui�P��P��P;L�$r�� �{�=�`Wp9��6��}��1ʬku%u=����i�Y�5E}��;�\ާ�l�����U@�͠�I�aiUH"L__a�T�h���O�+m�+�u]���G���]�`�T�~���͆z�+�����@S����I����O-�k�=�l�*�y	}9z�����Rwx�	ϔ�p����;�,p�����ȴ:Dx5����p��.�8jȾ{�͈ne����U9!�]6w�v��w��O������,i���:5}��c��uе�0���Z�䦝���	
._�$�M#{�1���� ��r��
mJE^+'n��e��8J�U���������<��3w����+�6{�-�������1cޱ��`��m����F���*, ]T+�:|����r=<c�Z�d{����v�w�)��)�p�tO������L�� t[=.�e�Ug���4"�O�
_��Ǆ���g�-h�|��F企Wk|z�w-��{O��s�X"7B��u`[�ө�i���;yw�A�Q��x2˩1��i�x��y_�T��}����d�f�B;[�a5��I_:H������e�6!ʖX�������҉N/�T������ �a�k[��|����UUK���b5kF�����c�~.���
a�������k@m�SF�=����3�̃9�Z|��^���e�=�e�/f�_��8Q�C��$_8��,K>/��E�ׂ�rX�J![����O}cui���x^���ˊw���W2�� �5�sC"�҆^�_6]�������g~,�x2L�@@l��}���D�c�9�r�({��[ڹК�x| e�??k��I�r��E@I*���S��p���*�]�=3
pA���&`���Q�k���u ��{)�+=/�-y��Z�)H�M�nY�[S#J�N��r�6���L�y�"43�%�YW"1�R<ؑ�Z�w�=f
C#d������ǦaE�uI�_�*LJm��y��TPP���N>����@�׈U^ֆ��<ae���j������ܢ�,���J���SZE�s��Dҥ
������������z�݋[i��^+uYW�A�n_v���>x�5_w��P-ܴ��p\��{6�)u���V�J�ˏ���{�*���F\GG+�A�Ą}QF�E&L`L���)k�Вe`�������ZhN@��5f>D3�6�q��
�1�MO�T�x�I<��_�],���rv�}W��cl�<;{g����]��1�ԁ��ḳ�.�џ6��֤�#�7gX�ODU�*k��ŨJ��Ԫ-�N5���{MZ��3��4	|<��m�d������%+;����<�w����4zwC�n�ㅗ�3�oF;�zd�E�RD�;i�y/[����1�:.���^�y�N�UO�$d.��>4�]7	�3U�.�.P�e�/QT/Ms�B��kwHƆ��R[���� ���\�w����&�:dEe��?�uD
9W�Ɋ�L�g/d+��(��O���[3.�W���x��ln�3�h�$L�xui�s9Y�%��[�H)ZNE����1UDW�?� sJ�HkI��䖣���ttg&��IۂڷX�Y�bi�WQӱ��Ώt�'�����;.���F����{��`��6|��*s��?3t��j����/��"v9��`*��%#�`�~S�p� �V��Ǹ��	�ֈ��|����$�T��=do�����ŪjK�w�\%n��{0�O�}M��31� ��Q���E)�-�V�j���.m�����ә쇚'^��P�U�.�k�N&#�v$I���@��3A�&�/�'��۞�kmaT)��a	ա��d��!�A0TȂ$xN6\����^�8�<3�aDF�;�I.d��Gm����`���@>2�zdpIL[�W����{Ìw���r�A�̎� ��}w?�0�/ᅖ�W��q70�|J��A��.�S��(�hX��L
��~�2b0ꤍ?��TG��ͯ;.�As��2r�,��DG�c^��-�;S�4?�d��G����{�m�9��M�GE��B��a���\�u�H�Vl��M'���]5݁����9��fc��E��ۮ�����Al�V�Y���ɟ��Vqy��Ji��
)#���]?d��)�mU��h\3�Go�R��ys��n2��*'��: ���(]�&������3�/��.���=�f�&*B��mE�T7�1��J	B?P-5���y�vv�3G����R�FF(�7��~͒��`��G���Ҵ�W�5�>[�H���Ƨ��p��2$[��u�ܨs�B�0�`+k�PP��A$���^�*�'��t|�,�B��o�;����z�Jצ;Y{Y���d���F�ˍs���dX�j�Ϗ�Q�r�@��_�l�t4����R��B�@��c�,P��؇q�d��]q�XJf(���D�P�d!f?h}��.E^r� ^�7x?T`cI���_���vɌ |	vC"℁E�'�e��-GH��~vK�M��ke���{�:h�h�IN%�d�/7������ܺ�|'�5Q��"e�9���2i0}G�����V�J�~�Ċ�����,����S��.{&E��G����}�T�0����z�2V
?M+sW�I������q*���­0�������^�L.�-��|r��)���SֿH/��ǽ�W����
4Z�{q!����oT�:��5�kw�5�|�h(�D^UO�HPw.Gm�^m�g�k�;f4�C�+�%��U��A�%Z��gA_3�"G0�w��y匈Z�L�3����3����%~��여?4L�@�H���H���6��^\��	��������(����kD-��.o�;��`Xk�јH��YS�)��+�/�g'�/��c�$Tg�5�rq�I}��.^Z�ғ:������YyD���Ƹc%;��1X�(��c�:Xt����V���!�݊�Z��
�+����M�y5u��ˎ�s0#qOE�9F�irْ�<�p�#ԗ��p ��}�i�Q$+�c��s���"M�i{�9[E���t*�#-���h�����뛸���k�3��Ñ/	 >7A"�x5ߓ���7�y�i
�����^U�Kܩ!9d���93!C?�X�K����'��Y�p�>�/���A2�=�풄4y��� �f�	�����PcE_�),A�ր����N��D�D&]Ľނr1��Pv�M�t����/[ ��@gRH~��S;��|�az��Ғ(��P��}y-"�X���,ʤ�������|�H�HMEP�P�"�[���;2�'�V�Y��&3�G#�?�T��>�d�ݸT(R��J�NG�tr����Wg��	=����b�W��������OZ��`v��cå��_��0����ȡ|�;�=��Zu��I�²r:}Zl$�0mFv��������1,
�� #�2��������0#�N{P�=�=R(���9r������|݁f!f�.i�i��oK�rǙ��)���]���I"�w���f��J�+�/�:[���6@�	z�=%�/ �����q�f�k��8e�����a�5�ds�w�
B v����D�Ap ����MAHFɛSS&7�����(�U� ���l*�ѽ=;*=%J%W'"No@��D��1�x(}�O��:s���V7'�M����ʎ�Q�s:���q�:����-�h�j��{����̟|($�����D����0�iC���HS␼���)ǦW�f�j�̐Ԙiu�����||�J����P�ET	����8��f~U��$b:�d\ ��_��9�UB$�_W��5X9�u���x�5�'Mmל(��U��\��)ڪa��Bf�:ڿ&��8:c�������V>��&> i�A#�(��R��Z�eh�G���D��zB$GS��5JP-	4g=U�G�v8d�4��
���%����ՎQ4,�.�1��Ԫ�p#+Y�P��O>����}yp���2̜ސ�z�ȏH�0�&��(� e�<�c�Z���9�����ݷ�ҫ�c�$Z�_���� ����1295`� �^*UU���/�`>E�G�Z�
g�6B�EM�~X���`Y�ng�`'ō�X���Z]������k�Þ���RJN/ J��)��W]�p���s�@���C*G�G�����E�z�ݽ�@��j���d�p+��oQ]�R'��: �����^+r�vQiGe@��j�H6C�L�"@��WFL�.톊��P
�6��
�'��,Pu����yZ�~�NN��!�_NK/�$�w�9�ؕO�d�����t�M�|���n�@�� �����x(�iӪS���A���?TȆ+��K�K/�FT����즅U���B�w�_��]��C�Q���{���m<x�YO������y��H��� Ӄt������6�}tC򷩻|�ZE���#�5�W�[uq�Mv�O{���V�&��#������>>��2���灜���{��1���S�jN0���R���O��3�:F"9`�y���2U0P�=�������h��q�S����YZ^߳�d'0.���(Pp��<��i.,���D���1�8�O���7�0���DO$j�O�-�`�[Gz�ߘ훾�̴���e�]]���jY�����UEe��?Z(��!=�h�Ƌ����L.r��e�Qm7c�\��/GX|��q�����)('��)g��Be��q�|��
���C%8};���/k��#L�0�fn�	Yz?�5W�}#�sF5�v�l��w�]�9݇�QKj��%=����b���T����2[�����<��˻;�_n�!����{a�H���Hp$�����p�Yh����Fz�eC��<���(�Hɦ�TNn��5k��KP����9{^�I׳�
>O�$�jD�y�O��:qT���PE��#�h�=۔�\�}b�B6���3�ۧ9��u)I`:#ޛtNc��GO`㚉�?���ݤ�Y]�|�Y�I�'��g��vWӶ3֔5�c�V�'��	'QV�P@�/V���-�q�{�#&;��Ձ���
t�Y��j�T-����*:3�s�b�"���r��^#�K��a��sh;��K#-ñ�]��s�yY����6��}"I�XC��[�9�E���~�횒�>9�$*��7A�?9�g�<��r��tw����Q;��-#�7.s)�YyFdR����>�є��8��ѯ_Q���/�VIu���p��E���(kHr�j-g��V�M�ʇ��C8�:\e��m,�S��{؏�	�>;F�����,F,O���w̝��ë���T^�u}~W��&~�ZQ�7+Y�_zo�Ò}�CS��"mT�&i0^WN��	�2z<���ӭ��gx=��}^�r]�ӎN�-��ӓ�T ��`�W��q�`���y����w
%*q����./Һʀ�+���xw�S�gp��Q>\®���c �a6B\yɷd�����N^�a|\�C�����(�Nb���7 'ܿ�J�e@kǃ �C?�y
`��x����K�p�no?�%����47("�N6�Lg[�l�R�c��㼬u�ў���>ô�!d��w~]n���
2v���[@�ˏj#��u ��	���^��7����"/K����:�}�O�Bpd.�=��$�a��(zU���N]�5�l���#�p|j��.l�0����t�%�o1{|��#x�����N5&�H��=[9�]���E��|<o9�J��|�"�}��B�6�@��g�&j��q��f�:y�^Ae35y,����6�Nu�I)�D�;ܷ�����7�n,��ne���Aӕ\X�V)[����k��)���<r��t�6���ih��,iՠ�Cd@�	�v��V�u��X�F�q�GMzT Y��oN�{ @���l0=���P��6= z> �/5�ԙ��!�Y�S�a�@�y��+��U\:[���V��=�� ���a�'+Y�a���Q]9�iz����)���� 3�[��j�N��fR��_��`u��4C�.I?Wے6	俽R���dݝUL���k�.��vG
i.T&�f�8��qh���-� �.��-�vv��"��U���,���2hX#�|2�J�zMZ&�Y��*YY�K�Y� Wȗy%���3|��X2�x�����ju�lF�(v]�����\��0	e�;P�"���N2��ں��h6�RU��&�s����`P�}��FU)3��\�yoT @($'��:C����Mv��u�s/a�]��̱�����¼Or�Þ@�(Git|B]�#��D?��N�#���Ň�$p�����-LT�v@�n������/9�~acx5�Q�I郏V��q��pmL�(�7 P�8Y����v�� p�����N��|���Jc���x�[`DO2��yO�l˄�<����ù��*7dJsi�u�ǈ���Y��?�U����L�+��┆�}6iYB�T�S�(�(y�0ZC�����U������(�9������F0�mG���K�I�P�3h����_A!�!��\���+�jI��d��U���D��!
���iA}i����N� ���~�Z����Mؑ7T�#Q����Ÿ�t��(	\�^�	W�v.
9.3�t�Ms�!���>Gu����V�Gv�N'Ւz��0��v��m#3L��)4`�����!�Y�A�e#*u����9T�R�)����`㩺��\���e��6ZM�[�˓���ɗ��<M���ğ�Ѥ���{>���f�h�X�b|5wdN
P�VH'���1|�NpRCT��?�،,��WO4����B����b�~`Ƌ���V1#u ��p���Bn��uAۘm�3��/W�\�E��c�����r�]�Z!-@f�3F��t�fG��2pF�QG���a�����k�1)���r|�xO!�PB�~��H�F��,xl^��+򈝑!Q�eCi3X��&�Du����d6GG���t���2UY%I���*����b���y���.4r]pq�~P���%�� �5g�}8�W��]��|$�.��C�=7��Z
�8���T�#4䩦���@�t�pb~�`��Q;�N�
�؆M��L�7�K,����M�/?#�)�̓)m�z�PAC���zVP]O�Iڦ"^\��Ļ6�Y�K�f��W��U�T`�GY��$�������ʟk��\�cS�.�e��g�t��
8�h3���+% �B	�&��s�k��$NA �Y� �\ٹ��@r�}bk��w��i�j���?�.C؈{��S�+�uy��W��nڐM�=������$�����!}>ll�N��Ѥ�n	��Kd�[��_��p{�[M�uo��{���QX�#�b�ڄ+�>�7��!�\��@o����]"�s���e���A7\��<�(X"�*�l�J�u���ë����t<���|^��m�qO��,�|��Pt��}ٛ��<'pP�~�,@"g���g�LQZI�Ļ���+���>�q&�炢�HJ�'z(\�D����po!D�i�ngv���)�V�����JU���)��n�W�	vb����$�F�p�p��i�!�	�`�[�&���I���/�7�7$��9L*����4���R
N_��}��r��iEt�*�9k�^���ʠ]���L1���d��`w�SN�d���`s�.ݲl@�[��
���Fl4��ׄ����E��s��]+Sc� Z�æ����������?
F��ڞ����n�˻-� y��l�
�r��,t~�L�U�V���H�2/sڃ	��L����.i=g�8�����BJ)��55�����<��n�.�a 8RH~L�t&}���l��).)�ib�<��0� �h$w Dة{p|�h��\���I,8|ʿ�c���[M�.խ��5�hl�#0��=R ˳2��v��2\ʨm'=�U(Et-y�ꮳ�rbڶ����l��6�����2*-٤XT�ܱ�\���~�����Ԁ~e~�z��OÜ���3]���2-���3:K��7�,�Z��e7y���]��l�4N�|t.HイڮV�^�?��4H�B�q�b.��U2>��GP��s;�Nc�7�89���K'���8�cl�L,��k���a�
g�,�&)���P�%����÷u�� 1��*�dx��Z�$�y�y�b�Z���r�U�U��r������y(���\��u�v�
�S��:N֌��^����}l<������1�����mi��� ����QԄ����%�y*!s;�WM�;��;pY��/n��:�H��x{J�ٻf'��ZB#���p��դj�~q��_&=Ω7�e�@�k(���H4�����gE�u���U�gZc��bKy��)���|,/"���3գm���JP��O����K�w��-�ˠ�c���3�^�mɿ�,�J����4Wn�N6�|�U�+��p�������H9>������g���C pxU$ל}�P�xM��<V�@����R�Si����A�z�7��6�i�<;��5L�ߥ�g���q&�����[[������FK��V�[M���
)��e^?�>�W��Ȝ,����=�Js�V'̈́�o�]���}T|�;��H�ߒ��4�N ��BS�(d����N��y]_��K	�
������(�+E�n�.�30q�Řk�%q���(���]�=�f�o�\�����Vb���=�y��k>[�Kz���$N��F��=*����y�s���85��vJ9�"i�{H��7�-+���dOw�f�UdG�*�z�M�h�-1W$I�t�B���D�b]���u��E���f�'+k�͸jP��������ro�Q�"Rl:�x��xb�k��i�>�[�R�\�xl^-0@�_4�$�W��aꥴ��{wM�~@�bŏ�����`\^�+_y����١;���٢�96B4��4�Q������<��b��
h���9mp��Jy�z�e��3���x�P[�t��@߲�-	�U���EwOۊ�!�+dP\�y����$]Ы\$މj�8����_
�s�M�N�:��_Ϥ��)W�rv]����ա1�Fs����]ƭ�U�S�+�r��+yg,�����Lu��G���J��(��뒿��ʱT��"�ކ��{����Vu�]�H��d�%u]ǲ6�Š�h����l<���g<�\���q6#Yw�O�>��d���QTh<���j�z�R�2�_��'�j�<g����
�H?�.�4˸NnW�	���sGmx��у��1r,Ag��O�����|F�6y��*��dL��w�?��`��a8�,L]%�/B�ϏgC7�U�~r}��\.1�;{C'?��; 4F�>S����>�?b�;߭�E��o;i��L-�z���M��f=:p� Vn��>ʩ>�o�{�K�Y��`{��N�O<�P5N f6��"���7H��|�����P�=/)p �	PVJ?�zd�\q����р:μc�4�.(�^��`RAc��BM8û�\/�a6�ձ(&��=(mգs\�����G���~w3�k���I���M�aIt{�3�&��;��hJ���S	�P[��h�T�Ô���%�������B��[���Β��UK�����t-�bÙO�\���0Q�2T#�
)-���q㳩�S�1y� �03�V���ߜ����z�s�b�'� �J@򇤜�=S��SG�әD\�V�6�0�=�o $?��)Dǡ��y��8xhs��ǲg���b�l1ȯ���i�⌀�?��	���}����{��g����������ߚd�0�=�Z�wl�t+^>젂F;����Nқ�lr����:�Zy4+mV[k��'���5Ax!h�j�h� 01"�0= j�׆���Wj���n��O���ʬ� a�M��rb��aOE���;�Rx���}D�D�gK����Y`�2�	�,�J�hb�Fw�=��M�ֆ�A�:S��}N8K�جl����5Ho�k�\��Ɏ��K�[}֒�\�qK� Aa4����)-��FB�<���4�<{vT�<�~�[}Q%�ņ�G�A�XW�T�@Q^a�|?���gƮu3d�����y�A�׺H�� �ը������X;̍�����W��!悲�;�L��$+�c?��5�o��/��,W�b�1`R�_�WC�JY�pR4�5Pf��о;��ɶ�5w����g�oy�%�)���<y��!G*,��R9Z�*�2
k8��ƫՋ?{� ���l=mǶ��
	��o��|JO�)
�M��_O� z�BH�z���݀��NX#Z��I��S|
A�4�4�`�������6����u�!��?���Zt��%�7���%K�u��*=�9MX���|�6ΐ��v%;ڈ��p�xڇ�|�q�\{w�\��S�&�q���j�rq:���3��=��Hζ���dO�B�|q��پr�`&dͅ�pt�I���~��-�7i� N�8�'G�Rŋ�f5�Z�2B4a�&a�sx�{B@�-Y���ra>��c���[��,�˚���(r��UZ� .[������[��gnV���V�2H�mE�Q*�tD��Ҁ9s�v��m��~?�-!�t��<|EEQP�Tb�HV�IBل`dM��� ��qE>��O��{�	�	U�P�Ie��00jg�aw������/P�ȣKկ4�7A�#ؽ�����=d<����k���Ol�����6љǕ�W����Rb���ɰ�Yz�A|�(�f��uo�Y}���H������ɮ�_����k*����v��z-Wv���&���2�v�J#{�4r�nM�bB|���r>����ƣߺ�0�9m�3e�h�lI;���ȅѭ��a��8=��@���7��-\�#��\w���k��h��l��_�_9�A�>�A��/�&aw�<����L����vpD��c>]�1�w�ۢ�d�����ְ��n�3��|uC�U�t�
s¾��HX�cu7g ���l�|Z^!||~z����v�!�6���V���냽n1�5i�J#c��[��cP�����5h�5[C�@ly>e�,l�"�ے}� rxTLAӒ�ޅy;���{y��+��I?�#2(1f�֨��:�unͰ{p�@���D��e���$R���X��5�;Mi�=�V��R��6$:F���}��%@p���>������d�?�,*�4*~c���������O�/�%S�x}����\��0��4� HC�m�^��X�T^������X�GO��U'�Q�e�9Ф����Gft!����]��xzA.1�&�တk�d+1;I~*Pu`��
k4��.\GwuD��Ǥ��tH����oR]b_{��+u�����f[[Rn�7ɏ`߻x�ҽ=%������כ�C~�S����2�b\��]��.�f�n�/�=N�PD�d	�:LS����;�?W�3b�˨HA��=�lv_��8�ڟNG+�;hV��*�M
U̿���L�:����P�X�:Rs\�<�X�]Ǘ�=,��!����@Y`�)�J�<��+5.�7|��xK�#��K�,�U���4q�ge�m��I�%刁�W#��b�'����YE������)����˶���&t �M���>A0~�_Ȁ/U��$M�ڐNG�ڮI٬`�w��c������|t.�o����mC���Cx(vr��f���B.6��F�w*K����f��:��­�P�q����1���q	ΚA�H8
K$ZQV�jD+��؏{�ݖ��pln�������J��bc/�7M�4Jf���)L��/*��B�WM��HH�e���z�E	���B�����o?9�ٓ��0��o��Z�-c�Xb+�j�Ո�G�у��������
�O�3��ǒ��1�!7J��ab��H�c(�/�P���]�]����=ߙ
�/WF��H		���9S�D�	4d��Km�c;sf��Ώ~8��l���a����qp���$U��T�AJ?	���%<J��*�tv�Ii����X�,���� �vy:u]��Z�nsM� ҕ	�I2�����e_������aw��y��=��\K��e�L
��񱦹�^�[����I|TX��2�4�b�	9S�dʅ�%��T�5ޓ;I�����N��ږT�6Cc'���8��P/{'�[U,R#&��5��z��`a��S�A�`<;��d�;6�p���Η������DqX��&*�W����e\3x/o:8	~J��$���ˌ�|��ި�r�]e5���1��[4��m@���w�6��K��k�'���#�$;%B��&֧�}���o �<V�u�uhrU�_�$��K�I�YP�`7|���ᑔey�����e�6��d���P���]x@�a��w/d�KGE�/�B�pU��s,�s�����H2�(�����,(���ϙ��
��v,&�k�P���;8�p���}��G�@��Q�Cx�p2p##��5Zզ�8��_&0h<#�n�"HY<����+�	%�p��s│��'d�'yʄ5C�(����R{��& (�@���Ɣ�q$M<���d}ز]��Kxw���:�I���l���c۰��������bJ�!|�,�%5���ѧ%��]#�����\����
��X�?-�g�ǉ�:��YsjUwPz��M��%?X2q0�r*���ƌWϘ��y:��nQ^.4�Rb�?J�.KDb�;��rl��}��-��������f�1n �5N�o�wR.{ ���to=@�E*,/]�hV#�ꂇ
����G��	u=����2�yE.L�O�*�8ڞ1��T��}ZJ��AөR���`�B�r�d.��0��vФ��v�4�N��[{�)��vX.���;�t)+���B��q� ��"����bA%=0K([i=�_�?�b�t�:]��۳��BH�W��DR��b�eP�`����ˊ��0s�ӵ����F���r��{r��l�у��U?����wM^��,�u�jU&En:)a�D�QN�l�T�sɘ��U^G,������+��e��\��ي	6��ь��Y7�c�{l�YX�EG;��Jꂎx��2��#�hr��,�v��$X�V^�g<��Q�h��r�/��H(���^dyx1b��c�g+`X�����h\��k���6�޴���#+��ہ<�ݨ��ZQ�L T����hW�y�An�Q ���ÒL�=����p���~�e�N�6l��_:8���(^~IL~�K��c�C��� �� �Mh���0V���F0��\���c����{��M:p-����\�Upo(:�1�	�x?PA�i1]fK/��lx��l9bD��$�M2q*d�e�șc�\xvф�!Wڅ&�X9��Z2f {k�� ��-l�Ƹ#a�K�P*K���-� ��xp?�u�[w�0�c�֨�Y�`�[>Zg{(GOL��p�WH�sЌF��F��<����5/vh �f�ӹ��I��Aq~�n�VՅ[�Vj���D׃L�Q��=d�@ܡk�7��]Pik�5��\(���V'\&�}x.���1�P[8 ��P�s�y}q�u���hL���Se�_D��ŵ��(�����fA^M/���aG;��~t@�Ŧ��֐��Y}�Rn�H��a]��%�p�q���-����`�Tz�|��m���혮�����gzmG�ظ;[tj�J��ѩ���z������5���kZD�r�ψGm?��>����G���ڝ���:��
G��m3��G� F:ffG��)Mj*߳Ao��)A��#��$Y�v�?	X��%%�R�U�{?���ؼd��>�f2����{�;����8m:r�D�#Z繠�����9Y�c6Eږ~e%z���A s�j	DZ �����1�\�e���h�X>�$�%���Vs�顨�p��d�	���B.
YǬۑ���t��J�>7�`@5gf��2���Eڍ�z�I&��s6rAӅD5��:�~��?Gwv�Q�1�|3?����`�7dZ����D�L�*�4�
M�OQ$k�5���)�L#\l�Gb��A'���a�RU� �j1�^�ןR�����.����?�#��5ڥ�l��ߙ���8��C�S� �;���;)��7�$�S3��t�>)��oJ0r��_JS?��L�-�h{�bPv��W���	��&y��L�����9�4>D)�(�j�C찹��r3����5�X���g�'B�h(��LPh�/�3w&����GQ� �����̓�i���[yEK�]8Dn�#��9"3nM%9�4��HtP%cx�:b;-w���^0�f]�vl7^��`rojTH�}�l��z{lq>��
�x����<�2{O�c �d��Θ�MvB�]U���p�}3N�!��?��ر�>"�̎��H3{�U�(b@�C��v#䎳,⺺� ��Zf!�UQ��5���q�ʰ���eJ%�q;��e7�{'	�šY	'��.�1'����{�H���������	�_N�2CB��D�W Xu�4ѐdÙ
,�#Z�A�r�ѥZ���7g�u"��!4T���N�W�S�Y^UcB&)g����	�ʻQ?���rv�}��v ,�K�� h�QLC�ǌ���Y�����I_�*"΅���l͡Fŏ��i���a�dq���:-!KW�Ӭ2��dj�+��;At�8�j��ϔ�b =w�Y�����wOY�5	E?Ϣ*,�K��.7>~gރ��Ŭ}��vo�ڜ���J+c����
�!�3�!]��5]�6����&��Ұ��Zm���ﳬ<��Kd�h;��ԁ�^9��M�~�D(�xA�\�|��u '_�ŝL0��\(��|,���`�߫j�jI�i������C�u��լdK����2�tt�U�<�s��#�5y[o{��r�2Y~h��N����9?�o��J��I����%�ǵ\`�X�	�і�Jy��a/�{!s:�>*�3�X���z(�iQj2�|dpΧ����t�\>���8=*�����<\<��]_l��d�jv�\]J3���'�֌m�d�ɭ���J�%I>c����*wȿ�C(�gD3O]��>I�Z1��u�}�x�����0��a���P�;W}W�9-�.�r���܏Ǡ��O�o&�&e'�'��O�e؈�Wc������.@4�lE��p���FehpM�4�6-ؔ���rXzD_�\�|.�iO��0�� ��gq��C;c�����[H�w��T��}�,)3��n�\�f���<֭�����Og@�O�%7���dn� W��=��� A�5�{����m,*/J�OѨ;�2��D{*�����Mg�%1n&�,���ۇ���tao��L5	%��L��C���剃G:)�[�|�3-�b<q�3���L�k;�M̩�.�ih�q��wVx�ŏ�G��������2I�L?���������yZ��r&����g�=c�KM#:Jlw����i�Ոg/sO�L\��3�X��
���_d^�R��t�QUS��)��h�Ɇڧ!K�����{�dlå0S��Ӆ���7�e3 ���?�R0��v�-�x��Q5.�]J#��j�l�2`�r���t �����,�����X�ӹ�.Cz
<�$�9�u+n+,G(�Hō�JI��� ���- F�C韧#׉CQ'w����ӥ=�L2�v�:��*�%�e�T	��^TC�9�� g���U�`8ω)����R|��V,��S��+�z�޷i��V� 9wz7���������;��F�����ceۄ�B������)���h�&���V�>=b�¡�R��v���[`c� �V�:(8��q�Y"�Eww�t(���j�xh�?	v��mCѫ���ڢyIE_5��)#���M���}W܏GQ��c5�Xcxh����F�]R��Us�G8��X����ёTx%۫r�	��J���5]B�Ɣ���"�s�@��Vx��{�ڏȪ�X�#\زID�w��.�=K؋�̧�QH9�{�����=lQ ��X�W�9���@U��SC�ئ��,�5@�9Zit��n�1	�Ҽ��y���N{B	���c�fw�B��U5Ŝ�3Q*Id8,���ܞ�a@5L�)�̑->ٖMXӗp�.��U?\<�'�~���G�o�&R[�)��6�o��N�Ge�fL� '(o�9 �!��T.��$˜���nʖ����#>�|��c�Z��G�" �B
�;H�i��H�,Eж�'16�F2H:�E�	��#:u��ʥg�P��KH�h�o4X|�&p�6� ���}���P���&Hɷ�`c{1�s���Y��Zy��,�;���D����K�ED�皮b�7��q/�1*���h����,8�+�n�;��)tE�U�@@�z��Z���F�q�><Zzb�;��HPs�$��/7���$��E3�Z+�Mb҆�H�5�%S<ov�{D�����&ᇈ�F@�[Y��po)
y���@���@ ���ꏲ$���q��C+�ct-X�,u	��	�ݽZѲ���gF���HW'6��8��-��Y����u�$�{��V������	�j;=rQE����?%Y|%�/�~2�~����X�kZ�[���v J�zd(<�����Ԗ|O��3�G�
�ZTv�q7��+�Ƅ�I!ثy�M)Kƈ�9��{>oYF�60���6���Ь�u�M�z�u�*F
Lu�j��/��RE�YYR%!��*�}�O�x��2���S�~���	˅�q��`�}D9H�H�-�aP{8���yicF�;����Y��˛�aVI�֩�;�[������J�u�c���Pd�~�iȞ�f{i����#@�];���~�gSKƩ |��l�u.�p4W�}I�O���	�<U�'�9��)����E&8�p�߸F�/��a$�LZ�m�}7���r�o)%�'6:KPT��5�ʁ��N�pF+�������XA�
*f\��}l�1v���G��^�4��p�R����ʿ�/6��P����V��Ԙ�0��у�e�Hv�Xͱ"���<ݬ�Δ�'�'i	u�~��+e���;��p����e�q�N�������{ޚ�v�Ҟ2D��:E�]��v'h�3=��t�0j#����W��?��՛��-���pj�Y���	�5�LZo$�UA?��o��e
���ݎ�U�m^ux6}��#��:�[�;q�L��]����as������c*�
�v]�I�9��+��O�mq؟�)s$��o_m��R���Z��jVB�&䄉��i#VwN���Ǐ�5��C��Ԡ��B
+T�xO�~;2r���ӣ��#QO�a֩��}�=��� �9�4�?[� {�ִu��1�o!��*͞�Ì�jG����|�Yf���Si$Ԇzv����8]c��2�Nq�&>� ]�.���w/�7���w�6>��,���yu֮p��(&��v��xW�#:�XI�ZAe�VkH|ʦ�4�»��y9Q�ń��s�d�d�o�¼"$�,D�<;�"f�znˀV.���-K�
	SA7���*��l�tN~����|D)���3w5>3�SIa��&ؙ��>��y]�H]��UnzfHġ�������	x<�b���Et&�i`��6����I�`��4��:��F"�o��R̊E*�q�y�j�I�+�H�'�֣�TX��D�H��'�ޠ��Җ�u�ѕ���,<+xc��vc\r��LT٬q�w���0�FӘRں�0GB���Ya,I�;�psH��G[\��u��7�L2�"��r.&��O�����:���*M�#C�C���G�܈0#�w������՚�d��0��~UF;p���vmܰ�Տ��[��)�q
	Y�h�م>�Tۭ�����J�j�-༢�c� W�J���4<qс��z���f��@�K�����e�p����ZM埾7Y��*�&�x{n��LI��9p���fd!��Q�S�Q�?���������*�Y/�%!�:�(w��I�kzfO���:x(g��uEO/R�C���G�b�_`f7ǧ?
5�L�&���.�zHW�_�ʤఠۯy(��=_J��\�`�ԟuo@3r���}3�S�	��J���;~�����JGj��GD�a�_X�����xO&��6����n�ZQٷ�n�/ d�&��Ӕ�Ɋ:��@��yϟ��_�yPm�oT�}�R���:��%�'I����@�fWD�#��[c_�*l�L��[�#��1�5��_k$�{�M}��4z����`�(=/"�� �	�9J܂�	Ob��`r���zइ�}(�|@��\�nFt����vss�2u�z�g(�H����Fī��4:�S��Bc��3'��E��t�f�k�L���%��X�x~��q&�"�Y�	�V�B-us,�k�D�ڭ�?��+���hM8�����|�`R��B��(;�rHd���=q.��2���(.��k��`#e����(��0ގc����~�y֋uE��8��&PL9u����`j�NQFu�53��v=40dy���-���_ܱ�>��/*��|�Ƭ+��Ϋz����vHѬu<�̓��'�Z�#]�W���^�-�e� o	�+fCմx�s���ȁ.j��9��!����� ;� F��n�/|~�i��F�?��a@;���K��,p|}VT���+���
eR��Γ_���B����i����\�yꊉ�=�$��)�u��O#I��V�$B�A��E�$��#e�� �
q��ޒK� � T3s"�i���rU�UM?���0��x[�+���M�q*�NC�)�zI����	s��(%�Hpю~��0��@lm��z�ܒx�4�<,�K�c �����=�;�Z��R�n��������D�NT�&�8̮e�	Ir?�����"�� �G��˜R�I�g���:ѫ>�s�B7���0q� ���ה�`0doYZє�8�bP�~�+��{�;�:F�C��;�X�?^��˔�Y;k���^�����=�����oz��xx�����-�n����ʞy��m�W;�yI\*�/R���o��ekGd��$��Y�n'�����{��<ED\�J>�$��'
��+�|+]|�-fKr��=z�z{0L�E'$��E���2Rg���	�	�~'[���_�Iyz#���^����ʌ�VN�Ѯ���0=�5����N�uί��F�l��)H-(z@�}��uU��[��f����E$J٘�����dI0P�O��@�����b��s{I�VЪ��L%Q�&>�8ɋuD2eBX�ŕ)����kx�y���X㔥�A��S3H��6I���!M���:�����
�ۆBӋ���LV_��K@]m6�VLr�w���3�{��=QX������[�Xp�D�Г�C|�X�]�S�<�^L~w���~�F�}���@���@ b&���}���D�c�D�BG�+;���@MB1z�_r� �N
�;��90h����ߎ�4Gw� 57@��S�*��5�օr��C@��� ~
�WQy��I:Uٶ�z����6��D5��YlP�;�&L� �[���_�I�ٝ�7Ы���ujJ.�@�."G����V��LLE��d� �cjUJ���#���l@	���xz�`��>�a�H:�E���CX��f��̘�P�B�0����z9�Q=ΌU����<e�l>��O~�1/�U�q#ITʎ�9��Y������MB�t��@���@�vvY�͟�=vY/Zח��yA۸��� u�:ւ�P���>�e�X��>�Ր3�ySf߽�k�ؽ�������j�~ZL|�]O!�SG6����&{�EW1L�;eƝb��4�m�1r��+Yy��d֪��)/��i�,����Jr�ю�;�T�=*������CP��5���D��-���j �ݗ� ف�oD�)w�@D���HD�i6J�%v�s�u�2�b��ӧ��X��L=]A��.	�{^�Y'�-���HQH%�Q Ii)?<�2�A%@��q���~f[U��ԭGA}�PD2^[�"� L�y�ǀ�0�<V����x+�@�E���� Q�+B.��Ez"D��x�
S&Ũ��&���~����5H'��4 �V��.έ�+��{�k��n'��WX@�Ѕ;�j�f�A���J�}fHU�n[���6������/��k� j-g�5xM,F������BZ���^`s�~3���6��
GL��5�"%>��]�����*����X �-��\�]%��OB�G�f`:R�.�8xz�<���/a֝����zA+�N���ďF2�r(޻+ӱ�Ʉ\��Wd��ҋi5�6�!>�H,�	>�Dx�6q�Q�(D	1疮z�Ӊ�Qq<S�0�(º�ǰ~���o�Tg`�q>���b�,�>��ǜ��-@+!f�m֍ fR�	Z�<77/<�k���-���r���y�@��L4���´5�B7�����F����9eѩ�i�l㇟�8��^����d�\���c�j��#�Z.�3�*���9�,�!e��a���lS�`�m�� 6� ܄�u-ua�|�sE_�&�ڛ_���������bC<�~�;�:^��1���������
���b���/���v� $K.<��=�@T&Z�Z�B.�&��X���48�M�V�s�㑭����AwI+�-\���%��`Z�Y�5c�Ku�@R�T��݁��Gsv<�+��' ��׿�E1���e�.at� [�+f�3�<SD��E�s}X�婅��6� �q[20����x���Xp6�M���l�5�0o����a2dZ��)*��hX�lsWVd����ov*?Qi�%|G>���R��޹K�������do�N�M��[8h G���*Z�[e$�1�X���$�\� ���@u�a1�Ci�E�3�wH(�MiF�2��d^44Z�X�B����P������<h�`��2��h�MS���Q�Ǟ�	խ�U#�*X)�*�\���C&P~%��&�rJY���*X��͢F֚:~�3�=����Tt��l�G��r��4 ���#*HW�O�^}��b�G�8�����t��,y���OZ��҄)�]�K+�s���W�����/ҕ�K��\?����ڦ�qJ��k�#�s�2Qu�����xJ�06B.��E���Jw�LS�&�ew]�3�]�s�dfr��.��-�T�]�k���Ӆ�������x���J,����ȯ��Vw��_�n��3�i���̇�.o���b��K����b� !~z��ݍ/�|6�F��.1�4����h����w�#8������&*ы�y��(�>����9������[&N~�k�Q����HH�!F�\�͒j��|&�rUK�D��������&�_�Fڅ�ॉ� ;�@o��3��5z����<��sMd�Ȋ��7�\����C��36�5xl��<�=j�4+J&��@�ǁb,?�׬�]7��=v�����G��h
d)��+k	Ng�H��\�ahr�HO2��M������EF5ja��uՍ]ׅ�q�vq곕��i��n+\8�z�u�Y��Ae���������{[�r�I��!i���hC���׍�e�w����Wա�s�:o��,R�����`/�~�$�#7�.�6���?:R#s�
��䞱����\۶�?��:73��m�7ˈ%d������wRHN�Qm�9�U4�������².c�r e���>�89A����̹ې�J�f^�h�ĺ�{/�?�t�%Xi��t�;Ul���a�zg�kfG�r�s'Ӥ8o�$����*�Å!tMY1ޢJ��G���b�o��P��y�k��~�e&��$�d�v� �]�y���l���:��to�Ք�D��� EۣÚ1"ُ!4�����^_�\�{f�Є,� ���-�Q���l�O��^��Vu:K�V��� 	��I�tD�-W̵ɡ����G�^؁���FE!�N�NwC��5�a2�N	���j�$��>����_���<M 
@�!u��pi�N����ڽ-�+l�ҿ{\09�O���RL�k�˛X����_����+��6�㜧k���i_�MB8�O#]�k֗�D�*c�s�w�OuA;���Õ:����k�%�����;��\���`���T��`�;-̐��BFy{ĵ��g�������dM�!���߲'�yO���iP��"!��`x�U�Y[q���c�ޚ�}�Ѧ��EUM4��[i�$�h��I� �v��"n#���nEΌ����a� )[4Yn�`���)f~B�]TX�^2��r�u6
�ۛ�I�Hmsi�߼����cc�����j�ίM�=��JK�Փ�r��^������-�iT���}_!K��T���-����	��X�L����Z���rqx\@�â;K�$��WE�V��H����K�I�'�f<�ÄVk\�xA8����$����a'+V���Y�����|9c�m��%����#�(��xW�n�[��܈il�{�Ŕo�s����@��p�c�ȯS�];����7y���H���'z=j�7k��Eޞ��Q/��������P�M�iܵ,��(f����q��1��M��K��*3����AnTY���PFE0HS�zV2��$j㍴M�5<(Pb�lo" f����i	0z��� љ���zZ��� ���U��)�5L�À���x]����&��kX;ԜL����gҁ'U��t�&!*v����=]Q���Wk2���
�Y�)N��ɋ�8�]�|�;�/�L�)�{mQ#ԅ{d��/f��w�S���k�L�i���z�6�>&�l�tdp1�u�tpD�yn�tv���� �偳����{۽��_U����7��\��������NM�FP�W���3W���pg�h��s�m�-�V�����}"���h�6� 0��g�0{D�X��)�):�\���sh^R��Z����}�� �f�T�f`#�e���k7��+V��)@�VA�wPRز���Ѳ�X'��w��]zk��Yv�O�������}��#���D��7!B��T��%����Q�
�c/'��S���S})k�R'�����e�+]%~��"����S��ǰ�(l�쫑���6�6-NͰR	��_%�\MI��:�{�0X�}'.{�l��:HLٶ�Ԥm�=I6��NބV�,KIk�L�"�����3u�{A�C�/�;��o�$��ys(�P��afE��xM��S'�m+�S1pvI?Z�5�`�~�t��s]�M��ɵ�J�t������IZ�߰]�ז1u��yU��E�\�x��.9�gX���=��`6�f�J�saE_?�Ƀ�_����p���^��L���"�LH���G6y����k�{tXe/��`{�xi�\-+H�X��*^G� �-��X��8�`��bޯ�r%�d�BF��pi0�0~騊J#��լ�=^�_�\r��>�w�5����ލG�h��b��(�$��l#WZj"��s W�m3Aͦ�6NnM��O?o�8�i�2�o���2Lh�Y��	�]\Y����v���_'\�!eQ�^�snIY�f^܀�ՍC�|�&���B�Z�,H����(D�[*��`��da,uzs�V�7��E5k�A��3�/�^����	�f+��L�(]���-���Iy�d���}"3��0�ݺ�4�DR�v��_�܎��d]F�!�HS|r��e:j1!����g������Uɜ�X����,C�Q�R�X��1�鞬���N?��gWy�6�܍�:t�=9[��b`aE�/$�ή�(�$ͻK|V����-�s ������	��UQ�A�hY#�y��cU���!W�`h'}��m���~ҫ7�s�z�OZ�JJ7mKu�����Z X4F�ʙftte
p���ix LÚ`�_(��[�|��.Ұ��d����JsQ��Ҥ(��'�]��n�����I�zZ�4$�3����:/���!�{�{Z���/�G/� ��h�G��H+`2�]�P��^]�1l�=�*AV���~6O#J��cX� _8�s��Aʲ�=.�/'����a�pg_��?߻\5sؘ;KCZ�_��)�i��I7�S��C�6ʟ|�$�.�� ���c��q����@eS4�� �<`��'����<�����jI��C�`N�α��}��`k�����,�i>&��'�n�[��L$��\d��
��KE{��.4� n4a�q�Ȯ|�4=�8�F�S��L
3�s���$J	�3��=�`@H��9ioYu�H���$(�-t��P���u�ti�}�s�Qqs~�P�^j��0��M<�<_9�j�ڊ�h�)�4�u����3l��.\'R+^o���6'֚���T�L�)bm���j�M�%�D�dկNK��+(�24sfaQ��&����o���3��#[�#ʩ����-������ܸm}�age��H��T}��������N
���w[SZ��6�@��݃vNJ�H1G.�,��x��[�yB��j/��/#�/r�Y���np���.d��ހ$�9�����v%/=�8�sOwV��*�it�+$d������?wR4��d{WKաS������#�4��룻��[��o&�vX�R`]�R���>��:�פ���W������(���-*��Ţ�"t �%]M�"��J���L6��¥�>��޽~�� ��J��ל����2��r@[���Xu"�#V��b��63�Q�i����C�WE!5�&G�U��[To%����8�jy�RutE��jAQ�<�|=��J�ѹ3�����Poy`���x�d�V��W�Ps�kz5_����w�OܡXH}p�-l�W�n�-�����&���ꉱ	
��_{"�?����)�Zc�o�����Ԉ�B0y����/����������dkUqEz��q4]� R���Kp��'�mV�b��y��I��eӘ�����- �>�NB[Y��f r�/��w�� �l��N���@#|Ԍ�E!�P��.�Y�Z�Q��$J���i$�?	-+$k1��1Q�h�y��z��Q�)`p0Dϣ��F�;�R�F�m�,�����Q��Ӥ�1�K�����9�ԍu�Wo��X�`&rE��L籮A�#�i��Q�-p��w��])/|�
\���d��0<�ZT�������S�Ϭ��ȴ�Q����a)H/���S��5��c�:e����)a�E�t��jo�j �}m���@G�K�D�b�M��?L_�b��2���''�<R�牬��m��+�̓{�@�DA��"R�����QI��@,�Y��z~D{M��㥎z@u�0W	�0������Y�ߤ!�
(��&h��x)0�#/������ܔ)�T�dB l�}���]�s�zU��9O QO��Q����	ȏ��,�q�|냔���t("1�{GG\���Mp���	)���TH��IJ�0]Y��x��g�#�J�S�s�t%ڽ�6d�\��jF!��O��vX��@$�խ�����y��K���O�hq
��s�[�D��
�Ip�:W���zn�u�sP�&���b�Oz2�(P����DK�/�^^�g��b{��\���*�@,f`̃����s�<��e�1Z��2�D�=z.r/�V'��5i��t��W��짂��>�y��y��ڲP�1黻���$ﱙLv��,�*P����hT)>�X�;��Q{�|����wq��r/n� � 83)j�	,RB��N�c�!þ\vG`�(1M^ViɝeE"�<(��z���H�H+.��?���t&�0�X���AK��
)� Ŗ�ͧ��"�X��V���l �4�#�M����a�T�U��|,�4%����OvF�[�e=����D��0�S�{^ɴU�L�#qRxz�(K=� 2�2ם�������)���4��Q�t�k��؂DS�`e:�������R��MD���]T�{�Ԕ@��]���'�V������HʍF��v�W&A��5��̔��d\���	��GVl�_l_��r
4�o7n���W�/iIn���Y�6(�?�ґ)��p��K�3����?�"���w�^|�9�MΉ[����C�|�?!�T��bP>���Ki�i-ݺI:fح�&g�I�UW��_RlX�9l�M	l�u�3�d�L������Ɛp�8K�s��S��A��@7�$�E�듺W�vv�Q�@��ws���r?h�Y�h�7P�s'�	�	��á싶���=�帊D�
�c״���"1���_�����]Gٽ֓}#Tx��|�V�u\T�8��q�9�<u�	�tǼ��$:rN֕O�[=˒���
���3Ž�k�;|
,�`㸝��QyΓ���RO���&XܢK��cג�W�ϮP_��]���<�1Ҏ_��r1�L�T]cqY��Vx��r�ۉ}߃Z���I�=U��[N����>/��H���@���h鸀����
�E�X�D؎��ԅ���=U��4��?��h�7�V�L��1�*��*�l&��Bj=�>��p�4E��0<߉��"Ԯ奜��[j9�cS�2��Z��8�H��D��.F5�"d��������
��\Y������q��ϵ��,���|��4��݌b�l0���D	���8{Y���#��u-�}��o?_s�$�#�6҉���<�����6��'8l|�3U��
	�zkW�S����$�$���j�����!(��51;_\��.�l����&S�CX���~<3$�E���<m����o �o���mB"Ƶ�k��e�a�������`'��g.I�3�����迢����v�G�0���������y�Vm-�*Sc����`nh�w�!��ہ�a�U�/b�5��$���i�ĄcNz�w\9L��Pԁ��ݹ4���X'�W�v��<����Z�P�k#�NY}-��z�#���B���%2~��OB��,�$���}vDU]�`!�<@���l���ծk%�o�i���L�-މ;���:Cm8���x���׾c�Q�+��M&���q����c��������l�N��,�N�5��yFa� W�����Q,*ڃΈ���?�.٦'J��6���W���|�9d�6��H�ؠ�u&�ze ��A�����S
�OI��1�m��k|o��HH�+;��lyN�C�F1�\����0�g�
W�����A��&0"`|�IP+�{� YǪ�/���4[̤�����qa�N��=�ߋun�� P�n�eQ����CIk�#��'x��&�)�ŊJ�f�u���٬h�K�ك��m��К�S����7��
W���������i+^oQթd��h�G<2L�!$�8:$Vy�A�nƣ�J��ba�n#��	���n� 2O�����A�:�����4�@�k����ߠ�����=��x�G�{�,-3����#s�߈���#�o��~��7��})̯)M&m�y5&��1��g|�ʨ%s	����{���b1Y��@�_M�7+x�aY�nh3�jD7�tQ����UT5�'
���vЍ��9:'�jXޚ&<� ����UJn\�w��8A���Rt�����[�P�t�%��z�ph�{�����᯷�/���Jx?�[5�r��4q�;�F�:�Qm JU����4k�FN%3���!�V&4-u��Q�8'���?B�M��Ϳ�{���D�;������.�o�\GMܗ8�e���S�+F��@Jn��#l��ʞ��K���<7,
�W�r�I�*d�z��j~�6;;q]UFE8n8�$2�i���"`2��"�"�m�H�qw�RNX�zG|���ꤲ���ˊ��8Ԛ�<��[��򨛅��L�K埾e��UFjTM�~���X�QI�:fh�W�kg��.��:{��0d+t��.��r�����g�uG+]"ɺp��!���������h
/��Cؐ�͔���tK1����f�a3�����.���,�O\���@!��e��e&i��;Ь+!��C�/@�כ.G�Z���Qb�O~���;����C��/bA{������7���5� A�/��@]���p=�
ܬl��'��~n�-G�]V��4�cX08b��f�4��i5��5F2VYծ|@��n����}�v�/=N�j��H.9$���^��MZ�Z}�T?2��%�1_��0T�%|E�ZN�����#Oв�6�.���O� �D+%�бwo�aDh��=0�:D��Æsh�?�	�FD<���ɝv5Ը�A���
��laO�
��Q�*�]��>�=�ə(c{���;��]E�����C�U{���`���hKo��3���@�ċa���Æ����,IWUC%_�+�R�U+BS�Ǟ���V)�l{i�N8��
@]pޔܺ S4�z���^�"ʝ$%n�2Z r|�M�I^��N_��T3.(� ��� �4=�E��?>�"yGSy�O�t^ �x�1�J�~h��#n�Z�ف�4�5��4?�(͞�=���x3uj��#��k�U��ٕ�&���-�УC8- �i�
���M09��0����`W��������(بi�K�'o��[&�!ڤ���m�ܡd�@�*"�H,��Ou VwA��\�ŀ`�g}(>�o=��H�����#%1K+�u��V�"�l��/�<�w����L>E�(�7���g��Y4g����������ǚ����U9Sm�+V�庫�H�ae�������q��[����Zp��ź� �|Q���c����S��8�ʷ�ڔ�ypлs���P5���9=ǪE#<m`�|�D�����X]�hp����v�e�.��+X��Y��-Om�O��YY��تHӆ�/��Uce,JaZl��a
��&�q7z���L¼Z�ӆ�_N�* ���[������lx���V(�ʥ��>Z��;ߊ;��H-.ę�Յ	��ˍY��?��I����?/�(H�6F�;�P6�a��B���?#.8�\�U�5:�_�a>�LuyUBzݬ��S��>��3eq����A���Lh�����ZAx>�oe�<lG�AX��e���_4�/�vD�Om_OE�"�L�Ⱦ�ML�(�}��.�p�F���Z Ϙ�h���}�K��lj^Bx��ʡnu`nߣ��h'/~�QS��[g�����xgW0+�X�n�k�w*��O����O�[*�i��X�AN��ӎ%����
a8g�f@��~���uo�Hs��C2�HɈޙi�M�x;����R����v06L�ɽ�{pT� .�
�=!�V�TO4��~QS?e����?D:Ng^�Ni��W3�8����7�ϖ"�M���� ��2,�L��r�������EJ�n
 (���ý:���Y<�@�f�����Yt���S��`0��U�66Y�����H�5p�D�/�H�*�CA ���֖/l*1��\:��yo5�!�9(��6E���D֤.P	�����ut<�b	}�f�Ǻj
�LR�凸���Np���.�/f�����$�=3��a%	Ư�"��@7��#+�2%~mPq�$�a����P�V����}%�~�s�?��J�����ͬ���˖y��̹��������ا���-�ϻl���4�f����y�L��a��y�~a���o����St��E���|�y�ƌ��_�T�,�����(K�+R����"�:��q�.%����P�?7%��f_nfe�&H%��ۉaQ_/�;��`H�A�,`Kc�D�(\B�8�@h�`��ś�Z%ʈ��#��kY�Gw���1L�>}6��N߹@es�$��l��k���c�ߠye�X��ӊl߀����T�%�To�K��v��S�U]��60@�������V|��Z����̩ۢ�^i�k��P�*�����]R8G�S���~^�0i����������4�@�3b��)(yy&y�H�e��p3�����aƗ�:/�mǅ�����hF\�w�)�0��C�g��΍(�v
��Sl�D�_�n����6�}Q~.��hRqo�%UW�`���0_ĸzj�A���A����4�o�u�&��/-�@y4��*�[�gO��Y�^t�8�W䫄�<���~:��� Iሯq4�rZ�"��uq��1�R���!^3���l��PK�五gm����\e�L�H�QPX���4dA*�\ue���dy>�jd+l�*=��虩�'�@x?D�U_ [F2�֍�	�Ӷ��&Y8 }
�����𪱿���;��~�� ��t\���Ȯ6�<�]C{c
Z@�c�:>��!��f{y��{�$�(��S�%�m�@b��vWZ������Q�l��f�vj��#�)��Q�ݨ��i������߼ʘwKs!�x#و����p5If"�q׸B�溈<e^_�F�`��.��±�k��+�Y bΨ��Qf�.�W�^���7m>y͒"N�H���G�i�V�tR���x� ������OG�^��|�t�t����ԃ���>X;����<��\� ���s�n�R!�%���
V�/vyB�v�A���p�z@\lm�Q��*Z�ݹ@�X��P���Ҍ�%��0a	-�(��t�G!P�B�,x�IC^ NV��Wӝ�I,] ۯD'��C�-'z,�Gr҇V�8������ݼ��Q��"�Ãb*�[��\hp/�P
������(^Ё)����ϑ�͡Z��>e^	��##	��$� ��fV��؈^�o�Ǡ\<4kâ�Z���9H����d���b�����L�5��aO@�À��$�ኔ�qTɎ�F'a�p�r�ȜR�!�G�z����Ѐ5ET�\H�n@\���J������z��(�$�P�{�k6����١�dۿ$�
��}�칊}U$΍G�)�!�� p}����*~z(I!�� ����bn޹zFL�(�t<̃&����?��y[��t
Q];��i˖��8��i�Ң? 
���cM����1QZ̷}�47��a�1, �aѯ�
C�ϖ�Na�0dρ
I��}�	��,%�\�������F:�W�j뚚�.����C��}�Np'�C�6��&r:g�޲��ɞ&�dFkr�Fu��k�lń��Y3
����-$.�%KIܵt�T}����1��$���le�?�� o�$�z���q['�����l�/'_"�
>'�N����ٮ�֦��N�=��'K��S~����s�{�&�M��r�_���+��/h�3g@?=��	�3�Z�}���'�!�����g;:�1k�!������_�=K�п��]��q"�n�3�:5-����R�)Nĥ��g���"0�=��
sڊ�8���d�[P,q��6��JB�z�ܛQ����j�O�'�s��L�S�H����v�?���l���O*��������<$ ����2��@��D��@��f������1�Y5�����ѝ�Zl�����L(|���sAcBl�������2YO�:�N0�j���b5�';k�nR<34�:�E���v�%�ڒ��c���As���"�ᨳaIݐ���r�B��[�~
N�^}cZ�$P��w��z߬0"�O@�nwb.\�:��;^�#�^��:�?�1�/S�Hb6�{�W<8��Ќ?�Jsk�NE��l/�n��\ؾ��!��A�*��!'�&[��¢,)!gR��d�dƌC:^��k�t�V��Ԥ�,�d��}�vl7X"�m��%��.F�\�ʯ>�wGۛ�%g�����VD��*�Z�t��v*Fw���V���kJ7*��T7r>'��M��D*�Z�l��G���Rx�@I�=m���a	������6�\#W�Q� -V�LW��^Nc���q S E`�a6-l��pl�
t�߿��=�+�r?��)̆��Q�5��U�)����c�8;��V��h-����ߨ�&+a/$tT��I�=&�ٻ��P����.Y�0l��$X�rp�Md'������MIV�P5IU)<dZ�i��u����drOR����v�7���Bfq)�3�L��|�-Ǎь��;��(}��'�$i8�XE˺�r�#�����������ZXGb���#��3G�!`�!T�ffw���b�^[��Mhn�����;�������u���vQ�|z�<�_��h�Y�.f��Q��Aݱ���a����k�ȟaia1��Wz��}�l�%tX@h��YM�b�[�X�+�`G�a%=��Pͱ�@h����� ��$��P?�`���}���7;���0�4�J��Tw��H�vxCGԞ���O	��M�''kgwW�,��v�(�a��s������8B�cO�P�Und�[E�9��ISY�梨���V3���-���6AEYq���WRa)���aU�]Ҭ����������p:=��R�#�F��/�>�-�����}7a]�&�>�(��xnw�O�YW#6si3Ռ_$l�Uxk����m�������IB��R[R��F���O���ܝ�׃7��bj���%0����6z�_ǚ��zb�I�g�����}i�6�����n�l���d��(�֜�j@�/=G8ŵ�Hq��$H؏^:�]t��,�$F->)��f��ˢ����I��x���Al��[!�~z�����-)S��Q�8
�M��x�o�%PL~���h�,�}�Ъ��V����:9���6����c/C��Q�:Ǜ3�MK�W���9�< (]�=��"�¸�Ɵ$��@AzG������A�UL�ͩ�SH���l�T�?�R_�Պ�4ꬬf��������`���faED2�j��1d�8��C��V�W�Y� �*a��znK�4�>sZ��]�`R�U-l�-A�,�o��T���d� �l(��� ��ߥ��y�o|��%�&��h�A}W�>\7���y�zwxP_9��P 4�D�<Aי@jn���7�R���L��i�7e	���`n7� xd4���q�6�O�E�{io�p#��z�x�?[]6k]��k�*g�8���FOd~�ʒ����b��ʁ<�ݠ��u��=����Bo��F�g�Fyͻ
��h~�d�Oq<�����b"ʢ�Ѕ�8�s�������ආ�\�"�Q�S>�r���MEԄ0�V��~�Q�y���&�7�����&�ѽ�Vz�Zu�L	�#�\C�nq�3��ia~'�;�1r6P]9�(��h-��/K�6�+��Ɉ�4�{6���D���U��o;yĲ���m$P-'7֍��
��}�8Wǰ�D�ㅲ��@#u˦����	1U�-tx%��b�)`}�p?c<��u-�wx����z�yw;�ֈP�pOo�W~�[o>�[�}&�V���)�%
���hɵğ�'�k1я^��QgRx&H���d���"�o��eK�7�bk"^����RSͪf��T��h����B\Rzb���2��l?��@�0C"���ů}Bf�/a�j�D��Ԯ�2���C�M�8��U�)U�F�c�UJ��7:#��;w�n��t�D�M��%B�� ض:�TI	�(�/���_j��h�GWQ(�nf�!�4��� B*�1]��i��Xsn?U��	|7���yVh���x�}�y�}���A���fd��>��9rŪ'c�χ"�
��#�#Oי�ڽ.�%R�ф�Ȼ����X��s;�G�:c�z}6����g�X����~�3�؛�2�qn�쭻{�����2��!a��w-L>M�~M��烸�l���5ү�$P��`y4��ZPEw��N9!�Mr�8ԀJk�D�]fL-8.�a��m�=$�����:�%��am�%Ѱ�ӎ/.nk���~�ZiO�h�J*�W֛'f[�Zu���{�;�kkڀ�y���i����SE�ɖ~F9��'`K��{�����G`G��_��J�^��I�y���t�l����<_o��	g�� ӈ�i?hU��gj�>^4�K�9"��!��E��fY��För �a}�BM2���J4etH�N*4mY<�OΒ���x��BB̭Y��G�^�q8)�:j7�f������Ng�nr�{.�ý�����<?��D	c+�˦���C��P&ȚM�/E�?��{NL�����">�}k��[��+���BL���=�F ��Ш���Dg�:p�X0�'W�[8Wz�r34H�2��#wn�������;=��$N�/����|v�f��}�� �3����GC�8�O�Lu�o^�Ȼ���f�%�K�#��8L�O�%5OPE�AGB.^�j�7h��Cy[�'Pe��J�����E"s���y��%}����vUfK�.'gY�� D7��6-^\[=���j)]Aa}�YlU|Q��ڻ�΢�����$�޿H�1Z1�6r�4k��7t�<��=�����E�<�����}@�&��q��/���a4��x��R��D|[;@�\�������EW�[Xȟ	ֻ�� �%O1ˀ3$H�� ӬA6��Ji/J����7HoVyr"�$\N-E+6�՟�/h`A/�o{C�=v�����mw ��|�j�w@R{�.O�ֱ��&Ӳ%��ǝ
� Xd]�Y�������i8sP������;�e��#��D�>G�W /y�$���W��K���^9���+z�&�BS; �-ۢ���CL}5�~���H#�sA�NX��3�"��\anH{�W�U@`1�y�_aM����y9���e5����JƊ�N~~�T�T���*����S�����Ǎ�C!d���#�� ����s�}p��]W�{�*~�d��I�J��C:�ٯ�K/�4����쨩��Ŀ4�"߁ߒ�Lr�+� �~~7$F�=S��9��u�� �Ɠ��dES�K�JWZ<tw�{g�P��1��B�<����-��:.��U�7��D}�(�^ڠr��Q@��{�K5g&����ߛ(�I>��E���-�a������;����̯�~��-��\��8
��W�T���|�a<��K�wuSTw��� �����T�
�x"���7���Kh�Z�2�q
�y���WQ67��GѮ�������,S1�|�y2گ��BIzU-�O4�*9��V<V��Ą�`ج��lnEȖfY]���!8bc8�uO���tAzĶk�c�v�R�l��L�.�Q��IO�,�P�6��R��f�v%%[�-a�FHQ����~��&�˳a�9ڔ{��Ab��ӷ"��n���]@`#KϪ��W�1�'a�i��t���� ����\u3{Q�Ö�X��	jN�R�8�r�)}cD(�m&*��������U��!*Y�|�k�qe�F[�$�U��z�������*��{Ui���Ӎg������:����;ݸF��+���jj/�䴴�w��Y�P">�^�U�@�"�+�
lx�d�Ͽ��&4:��W[GK���2=[�w�\7��8~=Y�م�����m熡��M��z�K�PP��.
��a�F�f7-y���h���̷[z�x��VKqn~,�t���J%څK�z�� �=љ�Q!��>�X�(�G���v>���hq��׳��)����8Jm�����އ�k(�hH͊R��N�Y5�A�&�2}Iַ��K��6���܅�^�P)62��r�h�m�G�Ӻ�z��0��&}4�ЙD�˕� �c�~\�$��`-���t���4A�
���fN�J��8�v�)�eDe�D卨�љ?�?俸�����5D�
����)7��[z��b��3�RtW�����,�熃#)�XX	c|<l��?����ZSȍU@A�_��G'C3(�]���k�X�:P�>��4�l��e��{�ОLB�KJ�:��%�/"��rZ�/?�c�"��0+���>��sm;�������a�!�'�>Y]��D�9ǁ�y��-�V�����x_���{�,���C��*�|�z$9�8��`���R��/ J3_��>���@C��ݩ-�wQ�'��d�K�ͭ�l��R$Y[a]��iv�9H�R�a8�[���ܡ�]���z1{�e+RȚ����X�xD�EM�J8����}�$�
�+�,ϋ��b9���蔀L|g+[ʡL��7������bƹ-s�#:Pcp\o���q>��@T��,(򋱘"���X�k��;!��n$JU��ց��������`cߗxR�,�ƫ\�Gˆ���%	�ۍȯ�}ط�j�Z~�e�3W���(b�q���<}d�bN��JN�F�p�������hو<�s�&I&
{��������)�v� b�m�KwʔUݩ�a9p��s�?��-������dn՚�h�ͮ��=��cr� �>/���E�L�	��%���莓
����S���-m�]��Q�O	��pYK������JWb)l��w������Yn��.�>`�uMQp�:��^����$,���ke�d������2���{�����t�A�C0�hj�_��2��U#����b�N�J>���#�{�1o}XgM�ׅzU�r$%�)Lv��4������L.��=��<b�%Ә~8�u��V,]�W5\��-�;Ї��Xݱ�Ƴ��r>�|��8[�˳҂�x4�~�g� ��({ϕ9��[���e�{�z���-�
�����H���0��'Q}���R���)`����������
��ּ��r����ih7;U�=�ii\X�dd��Pp������ǃ�cX�;\�.@Lg/�o�z{JDg�%�����J%�J,�O2�_w��G;�a�~���P+��a�Ƭ�%����6��Iz��ʧ����ь5��o�\�t��������zy����ɐ ܥ���-z��^zEX���zd5_���{���4A��d�$�ri�&U��M�d)�J���h�ܠ������o�����c#�I�X$���:ذuG�N����W�����p�"�9����1lb��ٖ8�jϫ!���:�׼$��kޜ<)�Vd��$~�!y�Y�C%!����@��յ$�:X�͔a|��F�!�+{�u��2F���e��f��DB�k���6�e ;�9��	�6=�I/�T�̰j�
{�7��#9�-MFrّ3A٤�Wd?���$�X�������$�F/~�ʜ�م� �
6�gt��q��O���ݿ~����9��F����[~L7�6�A�	��$�Ĝ�$D#\ȐD?�5�_��%��upZ���� ����^� ��a/�/�����H�$�id)��y<�"p!d]R����,7���e�V:�L�3Z����$H$q&E��(��`k3�8�j��+��nT+ơAh5����Q±�����/�
��5�w�)�S����Aű���P,% �wX���L����!����a�RQ;�{��ܐ��� y{���i��7�6�ᗌ2
��NpQ����Ax��&���(98'̆��H�M���Ė:Rob��Q�:��m��;��dh�&O�S���t���<r��ퟲ�.fe1E	�â���4�ҫ$�����	ͤ�/o�@1��ˊ�G͊�A �}����� ��sԫ��(�
0CwF
(���'I�J�R�$S�?�L0��qN�k҈�@�������9�k����URs@U:���!�b�yq�B��NӴl%<+Ш��>�$�%�AEr4^B��(�'7U�y`���E�Ue��ڇ���`�\�y�k�7Ơ���9F��6�g���gÚ~� K������!{ ['��8
����h({���e:�m<}]SELQ��M�%���c0H�Qs)���6A����J�6�M��&3vkiKJ`���0U�Ķp���֒���<l����M5*+�p�xⶦ��5��Br�y��zNx.�qi,=9;�*J�������}hd!
�]U�v�S�}a�"�{�m�@��"�Əb���Z�Z1�/������͉��(���V�O%�MMZ��w@��ԨR\tm�,�wf %���w�y�F�_���Ng��V�E�K�6˸,ʲ��6<�~a.-u����Q�Mf!������wy4�^W�7��A��p���-�n�`�<��rx'�5��5�q ѧ��I~Iir>����3��6~�A�o>�����G�dr��MT���%!��%���ɧ@�vh�x�޶T((z�|tS�����L@�cdvˏ�B'��!�-m�ƢY��Ged/q��0�e0��P����h��ۻ�#�%0���1�(8C�ۋ����,QJ3���s5ek�G��'ˇ��(�����̧��S&Va��/�g�9�Lt���g��$bT�Z��j__`�b]�խO�N���e\f/�����)G���t�|\��T��O��7�B�{����O�b���t�0A)y�6A�*bs�PJ�D�q�=ĥ��S��l��+�BFb\�UI(��,�0��o��H#-���T��X�f�����=IU)�7z���L��F�04���������[���xY��?|����=�N`��c���;���u$�f�]n����K�s�����	J��nV���J�a�{��t��
�e�5�U2��U�B�[���T�ա��X�>w`���mb�Te�{���ikt�4��z��K8��9 _8�"C��n."W�S5���P�=T�?�K����#�o�9U~F�M\���X��{!X �I@��~���'V���I�f���rۖ���6as-�&�������s>'��mY�*���1�� Z���|(�"6��s"������L'�U�Ͻ!}97o�X�F%+��D3Z&$�w�̥�I��
=��K�Fw�3�TL6˶<�P}��>��-��mO�oN��哿��c���������`����r�}����+���xt��&���1�������w�!��bd�{�TF��]=@(��ݦqo�f�Ѷ�#�8%�X�=�+{0TF����&g���<�d��N��E�^��Ȝc���b{z-a��	c�½x '�50��q��'}����!��6�Ҥ�\�'�t)�����$�:r���_�xc��wD<�3[	l��F&��1�&&O쭜'|�dѩ���{tɌJ���I�^�ū ����������� ˣ�F�k>�j�+.�!}/F i�:H��K �&/G*����Q���oE*e��g��O�쇍�S�8TR��(Wi���59�Ma��{��E�"��� ��ݘ���r�uAe=]'��f�?DQ�u�\om4?��H��O�S���d%/�~�2й��,ReKM	�-T�
��W=�!O�(����9�8��?���K��[Gztu���~ �,� �:1?,��`�	蛧ES�{��2�g_�O��g��kߜ����2�N�xA�a.�������?�i����x8?��s�v?ݵ;��.��!��Pi�����C�RZ5}Z����>�dz���R�|����j����A�d�s�+M��<�ԩ��'�Qs��9@:rA�h�Q@5#'(�Fh?�xS�;��V6��}4�D����uT��?e�'i"�v�=5���qK=τ�!er�w?���9�����vt8���BA���є~0�2�nU9��wtt�.A �B�Q|�0�S=8�.�a ��(�:��I	�@,G�Y�����'X�I�v�W`[��_��+��g!��N^�U���?9߅��j�XbԃJ�����V�N��8���% ��J7؆����P��2K,^�ɢ��v��<�l���ڜ3|ðW'��"����~jV�1���y�PD�ݍ�2Z*� ���߯�Z�}*�[)$���������3���{�+�T4["��c|�(O{���.ԗ?���웜q㑁�aR����擄Op-t\7}g�$��6"��A4���v
3U'��i���"n'Ղ�霞��~����'��l��GsY'��\�pD�K}�η,'����ѽ�S�IB�f���)�P�N�� fy����襼|�(�l{*�T���
w��v��EҳžB��r��~��Nd�/�w��k�B�	U�4�n���Ϟ�֟s�i���`#�׻������\o;Д�w��8��#U�cEa���z-[�^K�����E�ʪe�y7���'[�ܶ6���]_`���eE�$(��ۃ���^�[�2�|6c��%���%0�;ql��bJ�W�9��m�ު^�B��k��w�"��ֱp�.hqM��D�3�q�@��p_�6�Fd}�Ai]&�6�P!�p{d���P>q	^9[�0��È��B���w�}Ry��|(����MwVи�[�p�K� n�\<�����Ʉ�~��^�a�Ͻ��c�x:��]�ĉ�4RR��e
R����4�(���J�<�U]$dCCS|����nq�C�nW@�g<�\M�p�u%Ͻ�rE^{��í ����5�#|ӪcE���˓�Adt��5�-�1c  �.9)N7��:�~��T�SiD޼�3k�9誢��!�fח[?m�k��~� @�vn�:P:ĢY�&VՅ�]+ե�|%����_N��a��J�S�[����?��9����x��z����Y����{�߶ .NT�s^
5�(�< ��d�"���Њ˨�Z�J�-W�{���'C��a+Y%�4~���'��^���m��˂#�/�Y]�(쫃T�0s�O�dyGI`��GV:�?S1�J�Q��֚ۛt��7�_16��Bi���.��G��
z��㕠,��B��������;���yE\#f����#�t��-NW��B����1���/�3�S����A8���%���%��/��Ev�Y�ݻm���i�v����o���?�Þ���Y:k�^��4�}0�/Z}�C��\�Qd����@	O��û�3� �>Ir�Y�ΛZ� �ݧ�(mޑ2U~��x�E�HF��7&�Y16P���r�;�%Zw@����CE׷T�Y�t���;Hd�1oX�SK�o�B�o�״��8d.�=i���ϰ�k���ծ�Г>V��K)��Q9ܘ�.�=.�|ZN�DC,(��J�(7�Xúq�Rƕ���hK�<w~+�N9���B�������Q�qgB�9��;����%��Ѐ"�'ث���L@ʫu��G�m�c��$%ߌ"�߱�0��m{Z�_�p��e_�߽`�`�N5����O�	Ж�k7@.�@����eva�\���b�:�_���#��4?�H��x�W��$Xv�ĕ/q>��*�Gu�����/��~��0���s��"��B���A�8��4\z%�~���M�n��'���=$��5�Z��պ2�}���˅�{�O�f(T��MBH�1���5LŔ+�vG�*fx�_;����hM���V�15g0|\)�.��`����.�S)�X�� ��o�64���@g��=��ڎ^�{>���'��2�5��D'�m^�ϽN��!�
נ���Q��p%���[�pW���A�g��g��ĠaB��@����^&-G���` �%�*�+q�3�8��+�&%e��V��9��_�"@X�Q^
�AL6u�"$I�����ۈW����,����Ĭ�t�U)����,<H�$���B,��7
ũu��5�;pR `XE�T��i��5�&���3�ݧ������Q���.�QN?���9�W��)�5�bR�?�`q�M���j�u�`:��՛��m���A�ڲ�ߵ���cU�B0�o�ğ@��l�['��W��h�pG<f
��/:����
�,����B�;Rs��t>����]��^�tw���G�d�4p�NI�y_ML�A��L�L,�����¿u?���_��q*����w�'�~���>���+� �<���g�?�u�:����!=˕_��O��Q�!bF�i4�Pok�輯��] ��`#�$s��Y�zZ���2� HG�V���$�Ќ��̷s�I|r�m��l{��V5��lP�|u��#9Y�E<�&v]�̖삣D�d����u�;Մr&:g�n�J˭��6>���)%=�]�b2�$����q�����I��FA�2d��es8ǾS�CSw-�E��$����NC��*� $�]�=�t�oYg�N�5^G\����h0W�\j�A~�)���D�|���K�r(j��K�P/}�oʸp/�ۃi����qi�0sc�g� 3e`P׏1~����>��l�ƯҖ�bQ���b���7�Y86���7W�'���Mٗ���8�=�	�T�0/�T�LM�L��hp����?�?6h.�bK�:iN��������S ��I�-�nB�f�O��C�T3o��=� �aaa[���˚�Q�g���fFE���(���.lT��݊��T���C��r�(���g�G8|��;�X�!�P���:�"0�DP�:Ӥ���[{౲X"�F��oXW:(M��f��8�R���S�����I�U=���9�N�8�?Ɍ�tq.R�[Ղ־�dc16�\�Z,�\}�wE�bp�&�������WF�@����9����fHJt�.�&��~4:���=�����i��
�7n��;���M�D�W���`=�6�P �l��[{�pt�_V��T������B}�RBݛ��K�6��䏺�R�H��4��ǧ��Lt�*�
��,�A~�q)˵�A}VW%���x�Z�R]*]T����P6 !���l�|)@oupǮ�!�6��J���1��&���ޠjM���5�����D|$zG5U��6���Y�A����ۓc��&(Dw��6�@��6�k{6��"D%%�Z�X�����h��/6�YzV�e�^O�s��	�+�ہUa%���w��� ��؁���I�rY\�^iF�^as�y�� ������ ��;��Å�a�:)\л<��D���A�;A�=1���/�I *2�Ѳ/dܞa��D:*.

�������hog'=�e��ľ^�ʪ �Wr�XT_3e�ѵ0�+_�TRK��(6��F�b`�z4�2>�[)�q�b�q�$o��@�oP|�(U�d�<:���5ܔj��[M(ub{����4e@��.}y��/����l�{B���'8_��)���P4�~:�$���K��˥��.�5�}��$o(��E �0�ؗK����\ij%>�q��=
�Aż���P�OHe��`]�LR�FH��5`.�&�꿨�``h5��8z�duQ	�*��ȟ夾&G�uSg�_��ܴ?��l ����D#���A�ߗ>~���!"�`�⊑��->G�
���9ӊX�y�s�CF_��f���f�9j�w������L�V��j�u�]I݂Lp{X����d�����k�rxHM��[�+� ��Y�o޵���qM�ځ1	��jzɛ��S��.��D���<	���'�3U�b�+#wx�͠�:��c��%b��@�@�{$X.5&.��b�~� �t_(.�e$W��Լ�l�-0&N�b�|C�/�ҭ����G�q����Rgn+��$o>�x����ԗxT�X�q�f�a�Z+��0���� �м4�϶2v��M k���E^/1�/����w�ȊI9i46��w��SA͌��X=�{8���,Ք�Fa��?�1���U��`������P�����X�I�+χ.��O�p��J&��;6��ˌֶ=�p�ia&�E"�m�jQ!�t�	J��u�frICB9gMHF^��1��$���쐞l~�Dz���+Q+
g�n����mL5��7o]��>��W­��n&�]�7�S�=d5��?ܝ�����(����u����M�_o=�Y��a�~��8i�\"Q@/Q��}Щ�ȥo :9Cs#Uߒ��?����Q݉�<,�K�?��m4�.�ٮF�Xd�����N��{�$�j.fIN���ŷ�h��9=|���D�����R�\�I�J4�B�G��F��M�dm<1rR%�j�AMݔ��g2;��`��v3��R��}���G��9k0\B��J�'�
I���V可;�V��T���i�13z�������f-���N%U���s�����(5E�f���{^���Vמ�[E���,�#�e96Ո�Er������ߊPzת�X�^G����l�8�9�`LHA�8��&�g��	���Hv����7��,<�>�/<�"�*1�Y�7h�pi'Z�NzDF�d�WƐ�X���n*A�AX0�|���]GP^��RU߽���n���s�:��^��꒥-�s@�*�}L�U�!k{�2��/�ü�߮�[��/�O�ib,��jl��p�~��lq�*�y';�)$�������s��)\Ĭ�'6?��
bu�B8��ɌT�;�m�\�d��z��a~$z�݈�f֕��;����U�{�5���<���E=����0�b����U�uJZ�qT���G1�	����
�.�R�NZ{z���_�ED�mD�&1����i�$X���gpU*���l a�kn���Cڡx{-�=����a��W��k�{B^��|�Z�UȺ�?���j/��#��!U�Y���{֏��Wc�����:�7���z���)�����s!ܳR�{8����3��>�^8�R��	>{P7Q;n��#��s�{�\J�����Z�ǰ썘zYu`O�;'F'�p�(`!'��!�d+��Xؒ�"��e�zxvV[ڵ�����j��(���G��Ap3t�Q�y� M^�)݈�Qj#9�z�'lM��a��ǘғ/��ĞE���}\�uZ�M����ߧ����p���`V��>AT�ue؞��x���7I�݀�1ZΣ�~O��a�C8�lk��1�K`E���-�ery]�������T��0P����FSҩa�	!�����,�\wF��	�RGGP��e��W's>�v��D� �_	9�����!øC���	���N���r���LRz��TS�Lg˪�:\�>�_�ۤ�Ogw��1���9���[q�3H��$�\@L̹�Ʉ�}���9P�k#�٘s�����ү�ä���������y�1
�ܜ�A�����o34�t�c�X=�*��5n��y�Hi?�r���P��.2�K#QbO��L~��W�3�X���p����ø��[o�#����U�rq�3��"�n�@�d�G�&\/p�B�b���vb�a^ ˴��o�^��G�5��]j(f��u���*S��r�;�A�yQ�s�Z�՞��Вo^c=�cb�Yz}q��Y��.�b(�H��
���%!�
"���	u	Ӷbz�d, #��̈�32�;޻��9蹫�T>�nMEB�]3�E��5X��}p�X�yo-���0�Ň�/m	�{�jEe��" mz�Ņ�F��V!����ㇷ������ngH�&!	���>�j< �S�}��@iU�t�������
�x�3lH�k 2;k9���a�؟9b�/�p����.�#w�N;ذN-2ֳˬW���u�'���e�Hk,�))j#}�c4B۲�ia�D�sp�`"�
�&�_F!�G0	��G��ł�Z���ơ�nWo��!�gxe��/���T�Hǘ�r]�w��G�me( C�V,�ϝ�<v)�.:$+���4��k6�z@�o{g�I#3z�:*lje����R.Z��H릩�JVݣ�V�P �[�G�2{�*�����W�o�cE������@IY�v�O;{~����Q|�ky����j�h����ʺX�v�z���Q�Q�c����CE�ͭLB/!�\3�LV�M��/`y܌��\�xq��p����r�)�Cz�"�O!�=nZf�.Y��y�
�i���{5p�
���T|Ƈ]�<����N
�loE� ���y}�H6s�.�~�ܜ��5���1^-O�AS�h�3��dd\+*�z4��E/�� ��m0g��bk>c���Hvώ�*NT�Y��	�HuEtW�n|���Y�&^r��0U�o��m�~Zx�gB� ��d {�9�~F#P'�=�k��/o�E���� �b(��=	����E&4%b���0�Q"��מ$�*��r�);�>���z�E�u�\�F?]B"M����*��Z��L��챁6���� H$t�O�3z|h�~�'Æ������O��̭B�Ò�Tm��,А���I���V);t�Û�Ю�/�����zFE�RnA`�HHN��W��O��T��d%L���];����e�r�DW�U��@Ze�Y���oF��*�yy���K�)D���$H�wA�yџ�lH�x{�Lq��C��˯�ҕ�,�"�!�~���O˦J�[h�v�"��O:��z��-B��p�8���6Z���/�ٹǽE[���qTH�:c�_r��+�ݪ�C�62��h��4H<�/_�/Bn'�f��d�����n&���6���
����'pQ�MDd�bgh��F�&��9>4�`���G��ͱ�z�*����)�O�9�7&�@]=��=,Im2�2kω �/��������A/z���X�J�^݁:��IN�xQ;�Z� ?'t����9�ð��7�s��܎�τ#��&��������pk��A�����N��p��i�r���_l��4ـ����ʐ"�?��5�����#s�ʓ"m]�;�i�4�hN̥"�x�B4]�c>����0�Vrh��IM�C'����ih��$�Ѿ�*(9��׃�EP$td>�d��7��CTQ��)�;�A�e�m�Za���Yi�ܳ�ݽ:�<X�(xh�CF���W�ˋ<8'��:��k<����c��������d=@(韑"@5IƜT�i+|���0��d9�q�(�	�M[g���PJ�'HMe�h���ڿG��wH7��Z�+���~��"��/��c����L��h�Ru�ˣ&b!Y�5�����O��#�m�܂�6h8y�A�U�JmQz�������)=�����a%�zH��>.�#�@�����A�삉��N�61m�Q̞�_f��-8�Պ�:O�S�D��:2�Y ����	�cN�`�/1��(��.��ı�&�[�@g5��8P��[�L$�r��V��GN���|r�0+~u�t�5⥵J�(�}��6�+�G/|R�?_�as��܄ͼ�����ğ���~�����ɒ@��B����	��4��E\��P9����MI�]"{�BHf�T�yu���3��pz��Tk�<V5��ԙb��ZM�!�t0�a���ѫ��2�2�T���6����P��K�m*]�7Z�����_����dd0g8d��=�@�Hu@ �Zs&�g��(���L�`�Y�9M�s8@�Jv� ��oA�0��ܑ�pb6�wi�C����*J�nI��$��$���5<V�f��u{z�п�X(�=�@f�������^��`�-�̈́:;�����DHqH\}o���ˋvhZ�8�#�F�ƕ�}�(�뛢_y��Ga��E�����\ǀ6��&D��8��/�M�b��u��-z\(S��'�/���{�O �F���ND�=�?>g	nj�'�]f_���؋Kl9�[�1��eX��*�|�5��6��g|����	�^�q�HN�X��EW"�$+��Я�a���j>��75K�^���"�*Ø���|��+�ʈk���ֳ��A�V8s+�8�_�����mVj��I�Q���Ο�ѸcU�ݜ#�K�pg�2�أwW�|��'{�VS�s@�{
�S���ش��ڇnܧ�7MΞl���/ix�Q�^�I< ����!ˣk��7���[�q��쬶ǹ�/��s�_s�Q��Be\B�s#=�j�]e���|�ʄ:���%Е��GiI�;C�e�����������yr�=��}R�e`��Y�Z��c%{���&���m��f������d�����\F{.~���1JJ_~���eG�Z(a��uV}���vĬg�J*���k;֍��b�R����U�Z����䣞'�|pZ�'�*D�z��D��X߸ƍ��5/MN�{-��x�fˤ�_�"}azzF�`Hk���<	K�US�ob����#c��z��~q�kf����!�:(�᪛���B�{rl�:�,0 ��Sr7��(r+�	m���OO,!�4��qc�����
[���8=4؎'O�f�\��C�� /0����9���5��0��>�S��3�'qkAu*��	R-���oJl=�;�$�+�r�~Oe�j�V���b*02k=+���e� ��e�����X_۩:3a";:�>������ڬ>��Ti���:�;W8��ݥ���@��z��5��y�5����� l%�]!?���f�;��$I����o�S�T���:�Y/`��Um��pYX3���f�����짼������Jeo9(q�T�n��V�x]*���	�/�K�S���9�,��t�4�"P�:e���n��1��(eN�D̩~K����*�8}�Rk"]�Ss�JvY,�V�v����HDa��̴G�i�ڞ�ޟ�D���o�]��"�lC��$����"��li`h�"_䴬�����+K�&R�-5�^W'VpG���us�*3���9K��I,������^K&V��f�v�,?����(,�}��)9Fe�h�=����T�ْOVzCp')̓m �r������-��7!���ŵ��aѷ�!&�]��5▅���\��n+��7$ӌ�U�3�&C�	MA��ey���GkӖ3�����d��������gxY�z@2�T&�,�xu�������L�L"nϴ��7�i2xX�՘o3�d�����~�r)�e-��
/|��4�����IA�]�~��IA��h�u��e#݋U�T�V����=�s���m"����Ȧ�-:Y`S�M�5d�a��^�� �a=T�R�y�0�FR���|�N�����ǁ�� �g��:�6�� ��Y�u4C
	�M�5����;<؞��S8:��t	>��	4 $��>����#/L��z����:mYUߝ�a�4��:�OX��ʡbF�Ñ�*��Z�h��2ûѶq�û�M�/�	.z��I�c�%j��!��	?g��t���=���r+m���5��ա��m����a���m���pE������2B����i�<�#���7�e=g�n�@�O+j_��)���*�u��Gp�l�e�dg�������!)Z˃�&�N�"j�ې]i����
���'���$y�̥X�z���K{=I?��b��Bţ.u��z�E��$�D��>6 mҸ��2uP��E��%�c���k��%	hKU̿�V�r�j$7����[G������4�:����	^	�E���������}�Xʕ�Ir�h����Ge�q����.*������Á!�z�0IMf-[�Hwy�I�,�)��X|��(�A����h�qp$��"�a��M.�C�#.���.�Wk�%FT�;P%�A������5H�P�d3(^�Ѷ��DZ��$��x�cA���s ��ҷ����F%+�v�H)�>�fE�s�o8���Ԣw�]f������q��-H��S �$b��d��'�I�\��?N��A=�����;_���Gz��3�M��BK��e=�pg�4#t�?�Ȑ��t^y3B������T�y{)��?=�/��i�7�y�h�W���Ow0;M����*~����uqq^��Gk�ē��B�ʼ{*�!|%&k|\�1[=u�m����A�����T��Y��5_w� �c3�{��J s�edT�n2{���}*o��>)��muH�;;xq�ɕ��vY��^I_V���"�pq�u�A/�Y#�N�T4Vb;H��H;o�Vq)���!ڏ�b
��		�3�UFvO�������L�es�ܤn�9ӳbE��޺��P���u8�A���JuJ$�0��X���d��@�v�l�!]I����2?D���Y/���fr ��iהe:i�9��~e���]���
`@���;��>���U��-�G�(�uT !r�������]�ހ���ڣ)���Q\2�%����y���*k7�j�&[�n�yK��1j_P5�cQ����;�\�@�?0��<��g�7��<Ӂ�@��YK�����sC \b_�7
��4�"��%wɔu�=�ue�����Z>p�8����X��%���Z�����>r�J�x�$\���<��灑��\�ycP#M5S�7�L5��6}7܀���E#az��4��R�H�&�X\�Tz�~�r�O<�~��-'��׊B�P�������&��Ǡ��R"�?/�+
 ���߀V��*،eF�w�;^8
���l����X���d�kn��9�H�����`��nP�P��ȑ|XʁV�┸Y"��J����"���dG�u!�"�BH�Ɇ������&�(����1ck�h��`��05�R�^��٧��1���j:��	����.>�<Lh`��!���(l��V�S��Z}t#B���`2��r�~�jB���q;�7O0��K�)G�(�5α�>���ki�<S9��Q��l��'A�����h�BN�� h< �G�n|�"�\�]�]�|4�M�%��+9�Qo �R/Y����x&�R���c�[�Po�vV ܆X�6�5Ǌ3���,����|��'ѽ���袱g.[8S���lە���2s&4k%���%�{�Q,�HAK���
�y�p�tN�`�[\x��H�<���g'�<�~2�-��o���>4N���[�@��� ����L�0�������Va�Tc���W�@�N�Q��jX+)���}��Q���c��*"��#�ĵ��3�w.�q��-,"�t����guт\��I��C�	4�8#`�8�q,A�AQ�
#���-v��E��#s��CM�������!b��|u5	_@.�p
� ���M=�D0J��,U�_p��f ��!ZV��EX����mw���J2غ�'���ܟ�����p%#,z6����ц���� ������Z�6�#�M}�;��~��^���7�q��Őc��Q�=-��(gJ[_[��==	$rF(毇�����0���`U[���LfXm�8-�����4z ��ե]){�@)��n�qB��M��LM�W!|Q��x�]�|�~{ҽ}|��ʝ��X��}�.fHb|1������Bj�K!6{CGD�O	u�;B������,`�,�YU6)�n-M��*����淀�ʔ/����,��қ��]�)�}��4���j�o?b��k\{I	<�S���7J�,�A�x�������p���A6j�Z���g������ҡv>�H��B�z؝lR)�24�9�� yY�gm�w��8ƃ>�	,���
WPB���Gg�zU'��yZ�se��	(A�t#����ԅ9�A����ɖk}�H͓V��i@
)�!u���S8�x!�����皤��x���c;�N� z�B��@�Ĝ_N�h��`G��3#���cCaaV�(|�|qF��������8����wA�T�S�^d��zMИ���0���{���}�n�]�9����&��*?�Y���� #_���*�@N���&u�d�?ALwt��e�t���O^�/��2Y�9����&8Uz���m"I���H���|���{���ʴ�*z==;5Cg���?7zd������D�k1<��
��hm�E�A##��ѱDW��-�]�����BR�� X�ʮ�g�%����&����ZQ����ğ���a)jNn&f��,�%���8���N��[e���n^#.G�>��)�=�L��g��+��ӗz���4�eXe�I���/I
��p\��Z;���29fL2#�	��7���h��S4�h	�v�C>M�X����йg��+���~޲
&N��=F:��	�A];o�o��G�wn/D��[����绹��X��,~��r�O!��t���̨�R���m�FaG"�"�B� \~�⻊L+����"�������y	��-)d8�֗�����P<�t6��P~����L �8��NĕΧ��Of{7f��|b��]�*�_>��P�-h��$j ���Ǐ��%D���jͽ��G�#�����\.ٻO|��14�:愮Q��F)V n;�}��^ٿ'ŗ���f��Q��H��:j��X��ʂĖ@{~R�6��i���X#k�X�t�S�38+��?DYNb�28N�g�>�s&ֺ㔘J$�]���{���<��ǈەh&�@��?�P�V`w_w��mW��?t\�ꎁ���qY��Βh
��H �C�N�|??!�n���PB��u?h�z�u/��	��k���T���n�=v@��{`��ߕ5�[i����~�)[w�!N�~�ʁ6�Bٲ�����H�T�R�Uv��2��7�� [gǧG\/s�?�r����[b����-��W.��jV�far8r�n��
F����� *d�;=�2�K����b���j��5�-BG8���҄����	h� cR&�gLpm�nqO�c��8lO�׹j�����ſ`w��C�ߠ����/�J0G#�y�#B�s��dC���_X�蚞Z�7-ʁ��M��cG�+�?�^f�7����y[�D�*{�U�hRe<L�n/.$����3�<�x..P��h��ұX��g����e�
bYGX��0/Nm�Z�'�*y(���$j��Qu�����*z�@ۀ��a\��+R]�q,6�oD��%�WP0Lh���ɋ��/>�v�ƪ�i_��n��������y��P�6�VI�7ǰ��o>�=�KF��Ѿ0A��*AF[(�S���{�7a�xm3 J���I:��8�C(��_���%6�@��w��˨��M�a�X�6���T��E��s�%�]�q�:ba�[����4
X%go��Xr���4�tA#Voط���d���������$�I������4;���@F}B��
s&�u�gd�cC٥�'�
)��էn��0�{J-<�ޣ��:wQ+K�E�Qң��v�m�c�"���g6�YŖjj�4�'ځ������{j]�͊E8%�+�1��[����Β9q�iV��o�f���-X�D!�-��H�s��0�;�ҥJ��Ʉ�����j%���X�J���97��;_�K����	x���=���R~R�t��QI�c���3Hr6h)VXN�">�Q���~P(*@��t�g0׺�z�!w��d��R��t}��[u��ڠq����᫙��ʋx��+���% N"���X�Y�]�� �����X�[A4�PM*��D�2��������ޘ;�=\я�Ra�qJ3wǲ��[�`�QWs`db~�����c�f��W��z��V᝜ǰWC ����nW��YX�����O��@yF�a]K��rtd��4�	D����J��	��N���!5$�=#�c	�=� �T�p�}��IA��"F�[�x�[Kj�I�Aw"��;��mF���N�Y��c�X���C���8y���A�^�ܶ��M�/ox�_���w@mr<]�ym��Zw:�稿�\���,�>�^V*#Nם�p����u�B�)�,e0�A��}�w�=�Y&�'��!_|�}?�~���Dw�7w��)�h� ���4�6��X֥��!��_C��z�e�����78�D���2E�I=�?yu<ʄ��C
�����,��M�����2��#�Cw:�}�Z\!9�p$揇e�J�!]�]��:W����Ԓ�q�j@o�V�V���(��J����\�.j�KI��~��yhxK�JBJY�����,z����\�I?O=�����ʳ��/A]���9��Jك�/)]���={P������g����S�\�a(��c.<���ޢF��T9��K f&ƸP�LoP5�r5��t>��0Tد$��=�^Y)'���gc����*ttJ8Qrf�?/�X�3��I*�����9�?A��t�3�{�2�g��T��z�������t�3��� �pI��̓��f��ru����0m�M��no�;#E�;�A�Y��$���<�<�y�����ю$/�Ɨ��}��%�6��,ƕ���]�߾�p��J&'q%j��._������vv`[��n�g	��M��5J�L��~���j��*��yD?���i�iKO�����#��Jr���|El���������֤�y�)�� 'j� Ɗ��1�ci�,�4���:`���r��SyAV�Ͱ��� �mG�'��<H[}HS6w���qw~�O�5{�����
�4��ܘ�,^GV:~�x������wg��� l����c�Nܝ�6�6�J�L�Zc��w����)�~��\����8�z�,'o�yD>�efZ�/�Edlg����1�����}(z���"E���"��[�
�L��t'�E8�9��f��u� ���`X~��h+�Y��2�Q�#,X��bD�QH��)P���O�*!#�1�w?'��2[�GY�ƇRe�K�O�D.�_��[QC#�ل��:[�$��a��b�ō\3��_��r},��.I�.��H�%BI���GdT)��{�ÜjqCN6��X�0��dӊ"*⪫G��i�\Bȇ����V>z�\�T�V}Zm����@�6�Բ���d����Mg�l�h�2ϳMK�~@���;�X�Ox��$�d��&����2�z�ໍ�=IZډE~��߲r��b�q��i�h@6Uˣ���v"t�l�l���d�~�2��ݧ�s����.s��=�y*ӓ�ճ��ǋ��T�Y��2�_����|�^֞�g-K�ů�KC�0�RN�65i�a�)8wZ��p>J<Gռ` �V�M<C6"<t/��w���}b5���G��*+'���I��\bP��"4�lsݾ*ӽ��:q���aĵE8�Ş�}�0r	�6��v���yH������G)g}�F�8��Z���][�?���E���tI�F7. _�gy;�<x�Ex?��_8(�.�C�C¹B�G�G2��D����95�.;�V�K|d�����ɋ_`�����6�$d^ꖺ:E�.9T�������\�����!#��_��B�x�UO�׬�0�"Ǘ�֫�J�No�H`d�єc�,����R���$��DQn�.����� 
&�{��e�fA�g=ї7��5a���R�3bq�qM�3�+#pr��̣�]��f�$65�_ݲJQ8B��^덵
�x'���s-T�DE�1�0�p���������\�y�;*��5\�qlm�~*�Ʋ��eU������TA��e��J�M���AHrD�N��ᣒ��ܢ��p���-�ub�`�){�X@8��T�X��QH���RF6�����/��D)�)c�K�(:��N�f�1���%��[|��T$֐:��Ko���.�f��0x�wm���.��ˌFȞ�e�yA��Bn������/�Q-����l���`�m�܂6Vfth���G�H%�$�����tP0���Ծ%WBTxEN����__kk� �K���&��S{�X��̳�`�c���9�ɠ��/G�[
��ɉD/{@�Lm@f�į#��0�>�5�]�8��C4D�c���=K%fg7�3��ú�uه�M9��3���W�мl���p�ܢ���'k��w1��w�7X��^�H-��+pVD��7�h�Z�]��/B�,�Z{���N�Αp�Kn� ��n_\G�_q�9��/����yw�9�!�S�15]a_PZlؼU�{S�l3�*�R1��д�Þ��¬�����~π� ��f��m�4 	9�V����]����0y�ՙ�۲@�wUö�GN�6���c�׹����.�z��2}�3�R*����<l|v˺w��c��$�AR�M��	�
/�?n�B�89lzi�Ǎ�K��\�N��*vN�l����m�+pT��3Y�ĚĖW���T�FS\1��~����	�Pf�K��� �5�����j܏�����1�)�j�kQ/r�Em�A52f�&��A�"	�=B7��#k�FCS�������k[����C�3V�/5&�J�5��̵=$q�m��?����gMl%�W�z��P���ՙ�g�o���a��" �� �����\�+��Ůz�Q�*g��j�V��<KLMm0���, �:7�
�W�b�l����g�䥩b2Mdn5��n7maF��Z�A��1���A�ܥ��eU���S���ۀ>y�X���E��{��Z �����o~/��>��#1�^P%�y�ܿƽ"��@�5�v�j5׊�[B�����~<�Zw���h1��x��;2E�_�o&�*�I��:ż�sV�R��\ɥ��\ϔ���0h4�G��.T2U���+moG�R�S�Xt�Z���{9�8X��Y61����ʛp9��fmF\����dir\ʭg� y����N�j�9�i@C��麼0~�ڌ*J�k� p;���e`=$R�b)���J�,�<��C������o{�nm�o��i��[�J���>�8�)$S�'���wP�ø+B/��Ն�.���jx	7�D����#�_솘cF|=Fd�㻶�T�[�����w_^h"��Z$f3�zh]���(y���Y���� Fy�'���f�"��'_��-B�Sז�6��۸Z` �f�l2����,�E3S�@�����3ųGw��:�K�X�O�^���-g6W���Xs����k,f��hT��N�ae3��Br��+�cN.�k�s�J���"�ܕ;23	�!}��]��$ɧ��}f>Ύ�����FtsT2N ��[�p��ln%mT��h���]��/JY�����vLO�v��.����8��"��V�@�צ�C�>��&�܇���m�w�F��M�h�H��j�g�=~�v�*�����$�6�y�Xs�5���ƶ/~2զc"^	������G���IP��RtX tT��Ҷˢ�'_݃�,�q��W���Q�[0."kJ�lC�6��Uy�����Ҫ-�O;�y7�%�0`�Dz>������|�b6,�(��hL��՗
�+�4��!�Fa�-���=�k3bg�Yp£Yn�oz����)F��RJ=��''W�񂬠ѳdRx�4k�\2ub�vY��[������l��L=����doAni�Ny�qR��u/�6���݌M��s0+Q�o��B~�&N��杄Ley����V,��SH�jPF��c��d��mS_|~�d�N}J�R
�.�Q1-G`2����yZ/5 ���h���Ǩ6��N�9���f[� ��u�#h���|��5}DV���P���\�2�*]b�/L�V���ԳcZ�jZ
�}�e���j#5Q]��6=��2�jГי��V�{+��"�C�W�K�2�>KH�K���(ܚ�T�Q��R�y��v� �T	��Sg����e��dX�jLK~8v�A����z�y�.&i�vo;=4J�������i����pgw~��p�m}	��m^!�p3[�7d��9�O}��3 ��v�'%�l
��@,�PkPC�"�;	�c	�\��vGE�H��ɍ�rȃ���b�\v��뢫I�8���}B��y͠���&��?���m*�7�μ\P�}i^^1
�M���3�ǻ��h�Q�O��z0쪀�:��~�.(��-�p(<l��5�Ra��}c�E��m?�\��� �H/��~]AEu���A��t��?Bo ���B�Lz��}���{�Z��������f�U�k�vd�+���2����x���+��x��Xo�*��D��xO��u@���/�we����;��_�+I��W��ޛp�N�r�^DAH�>��@䌢���L�.�^�0�L0T���}�ܞq�$�ދ	1�����>���>�uh-&��X����H�F9�_��v'�ɇ��fT�!�Hٿ���V���UO�	"D�&��&��jX����L��d�ON�ִɬ�ު�/�0�i�k�����.��G�N���efw�:�� ���Z��ju%B�yc؏����d)Ӟh�\��A��
ÝT(���!� N��0Z�%b>��Dl����O׎�P�K���"3>�����>5�4�aX�B&ڜ?�қ/�4L����W�i�R$b��d�[��P����o��e��Vp��\�6�Q�)A�����0^4Dӣ/{�pa�e���!��`%(�4����s���.{ie�f۳�x,M�gFL�oR��C ��
�vu�u�wf?z�XFF�OE,�x� ���zl�Ù��x���V�aV8J��+2���Ê��H��j_PC����W�' n'�&�[_Z��
,�1G�����t��3�h4k'P��X�֦���0���S-F{�E��}�����+ fC�W�]�wgJN���ŉ"�϶���b"팭 �����H�'{����oE˵R��ec���f�.[ lގIU-�c!`��'=;��Á54���da����҉�n�O�w)FVQYkY�ҟq�k�`ǒ�*t"ep�ʳ��v9�?èr��5�U�ooq\jp{���e������XV�����`�9��Q�<z�tp��F�Xn`����
Cz���}
R:gDc�5�Z]������7t��~�;�櫹�ϒ�XF���v�+=��B�q�X�|�_$�1⤙�9]�0v��~�٪}Y�{�~m�>i�׌�]�?2tP���R���W}��>_��< ����:�af��6�p#�����[̰�7+=n��6c�J�8 {��\�ʕq3E 6�ߣzE���kޯ�ތ��2/yb��77� 2~͠
Y��8k8��=�i�{!��/���L�x�p���L���h� [)e"S|��>1���=U	jP	�C�}���Pb�ְ���$�N��E������1�������˴8ŀCC�|��q����yذ�c�����D��YK|��|��^�����A����>�@0��0�`��&K��v�ח����,��1���l}�>r�K��޲�˙�%1<S
f��l��H��|B��2-jX�~X�:�2��?2+[����p��t��(@q�Om@	)5�C�mZ�(�/I5�iL=mu�[�6�s&og��ܝ1��G�fDT	58K+��
m���s5�铑.���0�*��#N���^%�3�7�4��MD��[��l�}1��R�؁vB`����GU�����{H��z:żu�N��8��7�h�r�ە���P��//)D�U��<�2ѼkfٱsA9�Է��*�$�I������2���KJ�X��<���\�"����9_.m
�YwDQކߒ��ϱ��f�vk,MI��nW^O�>�u�٬�p�q�o�6���Uy��mS�x�㳘�� k{W�n��W^~Y䛙IM�BG�"�@P���Q $X�~[�'��*�$֤4�T	.�Z� ��S��۳����6�;�4#���j�YN��T�/_N����X� . �_d�PN��-�������WՕ���ty��w!^U��-���$��wt#i�*�״�߿�o��g�	]��a�R�T�h ��B�����~8�c�V��&ne��09�SsA�B0m��T,�/�4ɮ�� Ԣl���>�F�\;�F�p�7��(#x��pf/�S�J��,������)��²s2h�ˁ1�4&�a�����Y��T<�0c[?υ@��h$薢j�=�(by,�e�%<&;#J�sa��>��I~�P�$��b��"�h�G88����ɘT]��/�o����D�`݊�f.���!�_hv�`'x~�話�$@� ��:ȫ�����OB��T����J����^o�Wg��e�}E��7=�(�Q6�3�4Fx����n�WS���?�0��Ĳt�� �c��/�eom�<������I0ܺ�-�C^Q�錨x�N&-0o�R��j}�P ����F��eG�td�	�DW������Ӱm0B<|�4��c8�5�*���gkS|c'�i�<�����z,��CZ��i���~��yeGi��k~�R�5lF�0��������sX��|yJ��C�K>�x&^��O��0)H�haZ{Vi�3����kT��ٿ�$cH�(���w��D~i�z��U�4^V���f���dL�����C�<m�?�5���T����Zz�<�ҝ���K�KVpS��䋺�1ܒS�os�__�z��ɎQ�de�S��7}�É�<���� �I(�T��ow6�۩�
H�DlQ�ֈu@/i���3����s/��R�t�y�@,w�Z����<{Dڕ��ջ���ʨ{m���R ��`�8)m�L��S�V��-��D�t���}Nf+�� ��?���[*�
^#>�UR��=k��^(^4U��b�{�G����Bc<	���Y�%l�@&輫�C��ǎ]�N�J(v�{��E���RZ�)��2����3�wm�̥�^j��V`a�Q��=��"�.%C+�M_���b=PH�V�������0�]6���U�V��K���0Gu{/�
r䐼��cU#�݁�e�`��֧=%�4J��V�V�~�s�1�-���e��>�� ���m�a�!�t���f�j�XU2P����w8��Ozg5L9��G͏�]/�ߓ�¦����j�f@�_�W��W�i!�GB�cP���DIį`1ӊ����{�$t�5ω���}ڼ�# Zm��;�3_a� M�2/�ϕ�){˖x��{�j~����P���%��趶R����s�r륌uuyG��G͋HjHy��1��4Sۋ�p�k,��ա���
b6G���P\4ț!~9}�[=ݖ��AA-���K�2�^	��Cp�0)�m�#�_�'�d�'�q���h���1�����1�>�������K�E�@t�kGi��/�����Zj�Ӣx��f�o�
�����r�Z�2���"��a>���]��Xum��SR	׾��s�L��؞"`�i>�!s��P�I+NF�,�Y(���)�!�5��C?%�X�s�`�y����zj���A�!7���'/�"/[���-�J_uN�`Sw��Cݣ*���y?ϳ��C���Y!�x��UV��� ��/�&�"�u�ȕ��&��{q��[n8W�@f����s�=��7+Ӳ�N��Ԥ�b�P�_����yJeX-�K��F�F2D�7��C�a~�f�X8�9�s�ܩ�Ve�-��ULk��鮆�)/3�C���m㢴оS�g�bU8E���=��[3��YW����rK宬�|ej˧���O���x�e}��M�?�:l��-�{5/��d�CG7�`w ��ĥ����1v:/j%��K����M��f?b��t��~�'����{ �P����"�D7yG���v4F��W�����k���[��-ɧ����~�"��v����,���%add�L<t��He~>���!�|�Q�@H�����a�����1*�0�Ž�{")$�\�Cq��a��n�W�c�i���	u�������2D�A�0	�M����-�/h 0������l	�t���3�05���t 9�bvG?��^��Y8媾(��p�ſ�/Đ�����+TN����}PB!f��U���pN-��*O����� ��^�L�������&��~)E#_sm�j,K�k��.VM�Ĉ��s/s����n��!����s�&��%��f^Xяa�2�,O}A���Q�, �LcxL�c�n���� �G5B���Ck� ;�����=� Y��п���Y�cA��QzB_�gt�����X�o�C��~*�B����rN&��c(���>Lx�y����ލ�.�C��ǃFw����
�~d��O�U��,��xѣIp�r�#����9�6ض���=XG��!������[?���E���-~L�W4�er��7r�i�QJP��9
z*ΐ)�7���	���͞�������;���D�����^C\�^��y���<��ОJ����5|Hx7ځ �k����!���-2�}�^̫�#6�w)�Vr6.7�ș�c�/�8EAPt_},����tJF�~�)�m�ȴh�sn7P�~�l�'�
qfC"���p��8�1��ky4�4iz�s:��l����%�>�Bv���l$�:�6�zO�{nQ�ZEʺ�(_-�P?�lL�~^恼_�mnb!�	�L �#�?��@sI5�|��&�4��\$2F����M0�V��Rr��
7��YSd:�җKY�ghcK��~!�WiV�#W.��&��~�������{JS���l 4ao�ڭA��Ĵ[�V:���6�*=������dG��Q�<H"충��(���j��~�@��6�WD$�M,�����3���`�u�szO}����\�R]����d3�ۃzG☯�C�	}�y!4e�x����ɷ�v�5z6+���-G�P�(�V�85��W�4���)�l�}ޞ�O<l�8I��T�@C�r�{j� ������KU��J(�N�1��L��[��*[?�[�
��5I��o���06(W=��|k���*r�+�9c�b  LH|�͵���HH����d�������rX�'�.�z38
0D��낾�av��{������#�	��7���5�)S4��+��8�m��N�o�����O���AÞ���TX��A�����j��+2��B��X�_gcȣ<����͸h���k���Ì&G���`_�a��v���t��8�.�*��~ܾ��n�����%C��1�F�t��,uTW�caJ���tǳ-�D?Aӯ�m�:۞�`pB��j��J�[�<k��.ù��jxO�ըu��'��c�E')���]���W��DS`1��J��hp�����JD�9�kUB�� *#����&ڕ���:�wzt�E�oV�/����.��R����W�0�ӑ#�G��@}A�T(9ګ�)���Y빺�O�5-^���苴l;@yh�\��n��Dщ�N�M'h�Ӭ����F
GՆ���=�O��춁���ɉ̡�RT�I��y+GP�%�d��o�w���[iuW.�%��0��>���8�?<��tc���`i�V�l�L�`�EM�߇��1Xt0�q��δ��bQn��BJF4��z~5c��#���ť��	�]-�������b�$�!P�q��Ǩ���)�9�&��F��,(�m?�ï�u����j9�!���ZCՇ�1v{����T_�!̱x˸`���;G��Bܕ���40���������S2SY8�b�\�%圵��&|�-D;G��I1�����o���	{S��0}࿴ԗ!(G��T��U��uu�k��g�gi�* 1���J[3^ٞ�uԌ�4Һ����
�z6T%�2EeK_�$�|F*�XD@�L����:��#x�DQ�Pm���"8#����LO-��%+���� W���_z�,qZ��Fǟ?k�Ń*o7ox���Ήe�!��΁ǅ+�{y���P<�4����G��v���eS�K�^���[��3�L�,�@$�M	��!I|D�	��0 W��9ZΌ��B�J���Z�y���5������W�z�t�܂��g	~�����r�/���������M̨��l[Ҝy�4��>������
P�SY���Q
&���0�.��[�	�ד���ʹ�O�`���9E奖k)�NXm� ��� ��<Y�yf�}p����k��1E��^,���A
e��&�gTO)�X��3�iM#�;:l���@�V�d\�e&M�5���=�e�7~����h�t�^bS�T���Z#'�^��ŵjƠ�ut����וb��4b�; �,�oI�&�`D����f[�n���I����,ͩb7��� h�@7�>�;-�V3X�.�-�/�?��$�/6����!�K�Hsw&9����@�j�P��P� T �����B埤3�,�;j������96�T|� ڻ"@�S)�{��8!�<���JiE4S��`_<��:��S�K,���!qr�6���qY��� �b�VU��Ә�� .�?�e�� �Gm��;��l��Cfka�ڰ:��b�0�{�/�����-(]��C.N����J��C`P�cY�̼գړ�^������-.�Z�$��� D9N2�	iY<G;��ٮ]N!�I�x¢���8��g5Nkx�mΓw@�&��	�f� '�h.�^ǟ���-͵W��������?��D6�� qQ���obK'3���O]%c |�]���諴GQ`���Z��y�;�9������7���8�^:
����e�]���d�C�L��c�N+��T,�q�iP�M#��a/��qW�<�n�ܧWU�S1�3$�w�K-��iv|��db(�s
ނ)��K�T@���ա����=X������!��!,,�4��+|9o����UV[~kᇓׁ���)(<�����&.F���6�ӋF����C��m�fzy�U{%�f���n���'
U=��5M���=ƭɘ�Ɇ�Z�ѨB�x���5ք��������Ū~�Hr�r#���<��!f`�v�YOdu$�
����otEՅS���M�N�&5�i��Τ|�������0���1��9A�	������t�tIZ���a�8Eؿ��Z���7T?��r����./~���K�$��Dl�v�;���Q3�w'\"Y�{L�SI�Ԥ�ꃨ�e�<Kt�v`����=Q����.N��p3[#4W��j�W�4Mn��@�hK�"�%��l�����qX��,�����B��Xw �L�V�"b����w��m5l{�V�$�jE$�rֈ&dA@�a0���_OjԷ�J�x_��W�'<b�i�%����W�*>�g��4�c�ûhH�0u^v)�~-;[ƝF���D?Yge�b8+9�c���	��<�o�H��f^"	Ձ��8_�$�r���^w����i�O��ʭ�J:q,^"�ڐ�_�Q{w2�pg��2_d��|��� [7掖X�����J��'&r[���f=�C�l�H[}f�2ڏRܜ=v���73Ã���l���w�����r��U��l>lW[(��զ���B1J����@)r_A��^��]׊^�����\��ZQ��ւ�t�����>)5��WͰ~�w����:���բA;����&hp4-�G�('&�#�#�}�{<R�ʕ(��+����;��:�q0�n+~��V�HF/���_8%��|�����V�V��37D�u���o� U@Dy0�[��G�'�񹍢�b� � lu�+��j
�J�i��o���1�X��V�o2SQ0&Vz����bQl@�Č�=.xv�R_�z�K�JcE��$��*ڄv(�gw�%N"14?z�3}��XV��ǚ�u�5��!'�I���LԮ�X�T���o�5.�j�`Sؼ����#}W�����V#kп��	�}�� ��W��Dv ���׭�TAϤl��Q.�,�3+�AmB�B��I=��z��[��h�hN�~��b�J{��0��K�R�T?�@��«�Z�����봝�}c�ꙮ���<�Xv��p;EF>#2pv�ݟ;�b�xNy��m��,��HpeѨ�k�T�`'&����J_d�QG����N��x!7�]�=�����r�){�����r�Aa:=�[(Np*π���N��߼�~�&CA��mQ��L���Ͷ#aF�&vK�P\�DnBc��r�j+h�3A�y5m��������ƍ��[*����)Os���+V<�c�t���U��oc,A/P�k��C4�Kڑ�]_�JO$����oK\��ְ�1l�ť��vs�Ԛ�S6�`]N��p}�/��N�
A[�'��;�gb�E���p�}?��e����A��=�4h�1Pl?��F0�in��!-j�p��*����`�P�й�� w\'F�n����i<)�N��e ���'E`�b,N��~�XzC���a�E�;b
�� d��E��9��$�싻w�\t�5'��c�/<ą��O�_L��y�)�an�N|0 sS�����[>(1�����*�AbzT��YKXIK)d�g����[ö�r�'0��&"Dz�E��K��DZ(z���1�g��@��ar1���G|7MF{���^�C'�(��;1�E�<>����P>�ˇ�6E�5g�fB�(q<�3e�O�9p~|K�̘s l��ǍQp[�~e _٣b̮~��#�|�a�s�C5o�Z��Yg�鈘?�	P���UV���Ŵkw{�������F�3��S[㾪)q�4sX$�j�rv[���`S������TR�K�٨�q�&d{!���G���v�7BN��ٱH<��?|��~���k�%u�|`Ý�+�r)ƹfz�H ו���W�i�Y��0+y�^}����t���'��)��z����O�����֛�cHk��$hK@
j���̙�:
�A`Nc@
ްɫ~v���BяY*���-� �j%�{�B�i�}����ݽ߬K`���g��Ҫ�80�<���iQ_<b��6�7�� ���6;X��h({8�C��n��r���c�X[3Jm���*0V�K�n��H��@�qnC�e*�E;(4j�B�5p]�*xy�E�%���C~�Lq�t%�8|ɳՃ�Z�m�.%�!�����`㯏�,��������L0�\a�B�T*�ς���y?���1�%ꫮ��:��О��~��u�����b����s16����EĢ!^g .F����~���c�:l��*��c�~;`)m��8H���F@�(EN`U<�,2�1 �c{v8<C�Op�6����^*�����<#3�����GM�֦\i�F�b���0t�ի�;�nI$G/ˉ��i�y�	�E�\+�w���0X��Μ�r�.QN���	W�z�adrna�ګ:g@0��)p0����	׶'����ˠ���5޵86x���R<Us� N)�$��"vn3~���p���x?>��+�\hj�?Z�n���l|iY%�Mcz��N-��ܵ��۴�J�`�D�<����=��!��H.cHp�$5�w�]���WI�}V{<lG>���G�a�Lo��J�}�Ȓ�&
3fS�'k&��?t�.l�1%�l{����̨�?�ܐ2ov�l�s��aMH4��ʠ}��P���A|���%��]*hJ[0mdj��ЩXh���$���F�o�X�8�o<��L�jRi��z���=��-��
�Ş�yG�A���i�~w%���	��;N^;�S8��˪��L�.���Ѵ۫�\s��Ӫ��{����t�BJU|�v6Kr}�q���6bk@{��o)��O|�Ea�X�Yצ�D�+)��ȥ��%�|�m��ux�U�:�T�T8]��@�wQ�ON��؇�A�	nu'ՠ�*��*�ʅ9i�W6�}^ߚ0#�� $�Я�X�<���p��^��b5�RvE�� jT�E%ޕ�QV\Bg��o�r)�9&<�ՠv�A<4��2#j̼��\c�&�{��9�|��i"��~����]�G�Ʊ[�􌠃gوo��dmL��.�.�~�9hQV��+¥����%3p�� ��ی��͜j'�te%H�����.�)6x��-�aA���R5*MXV�������X�;n�=8�V��(��V0���9���]Q�p�v]IMKvA�)Ky��Pc;������'${,�����<��c�k[B���*����/�wh�G���r��*AnC��ե�ѓ�UGR<D� Tk^�R)̽���yR�aA�ѶmL׏-~�!������~��,6��/�*�s
=x���]mmt/Z�S�J������_1S�1�;fJK�5��Nv�3�zs���0=�od��aM�H"�[d_P�]�Y������Z����9B�Pm�~+�"��hd�����T��ܙ�U9�Қص�X�����g�u��lm�ƿ���.��J���a�?��et�Lz`uLAy�N����d��,'�����$��Cȍ�^*��.6�4U0݄����B�.j����N���w<´����f!�~�\��$_k�t��=��.��->B�z�i�t�K�
˾��9����c���I�ݴ�T�#����,��6�(�n=}vp����l��V�ɷj�r�H�[,#7����3�}:(�(z^��#���̉�vtDVy5E6�~0ů����������z�������(t�����k�c��{=�J�� �*�f�Np�)}_�N@������~������\à�����m�`�{�I�*F}����w�7�I�&�0�b_�����L��ҡ���z�u��a6����^���]���K&�9���omқ��{,1u�3�2v�p�;�R6(3/�xtVԼ\���#4���u��� U
�Q8�ʌM��V춷f��|Tϩ�_��`�e����P���yx>P�p���Ԁ�hk-���,�m�*,�x�g.����X�X,z�c;�y����hDx�K�Bm��|�d}P{����0�L���փ��M3�v09���k�yۖQ���57�P̱�?l-���e@0[g�U�%���Utt�����r�2Mر���~��~���
k���0��>r�J�pw����\]�ؠ!��>���)Z2R������o�T4>)/Gp�.�,�����}��nW0¦���T�����NB��MO����"�0��D��n�!��Z���Xj���"x|f��=[:�FT��7lEvx�m�i��A����K|b�8ݻ��1K �{�v��2h�Hb����������X���4���*0x�3J�b)��^�K�|fs�#"2��{�$�.}�{\�m������+�aB"���>ۢ<��(8�.�D�̋���� S���2�[_��:YL=�g:����3偵�W�H>����$��9G��ܲ:$|A����ء� f�(x�����[DW���;�W_�in3�,j����0���}���"]���_�^f������Y3���1Krp����͹%_ y�яK�>c 	��r�F�!�璡�KiZ���v�/N`ʿ�B*�>F>	^�|L&ku���κ�e������8+�欇���.�Ā.-�wŊ ��0筤����U0Q�F�Zm�UNܻB�4��Jз���b�F7���#o�/��<>���|�ւ���UU��,�������I�ef_������c�~��Q{�l,\�4׸~b����v3U6���m�(Ϻ^Ѷ�t�h�SU��gٖ�m�m��5����Pеwp����N�� ����u#�@��3��^S��SZ������r!� �>$�ж>�R��h�2�G��.QO�vq^C�����,'R�?&;���"��޶J��>b�SNdt+��W�}�|�>WiO���̓�w���Yq����j��J+� ��%���,i�`b��b�άA�\�����z�G�#�g]��Mb�>l�鉈�%e�ǎ-E�=��"�#Y��H�)�	�١�j�8��m\9����q ���!'F��4I9/��=11v���������!Y��M��me�0���W���1���V_}��|}��j����J5l�t��]Cm����b�4u����a�~��K�#�T��ܭc3e?��*��M^���xM����
���~�!'�Cﶀ-8���C'�f#K�Ǭ�wj"G���إ�m%�� �3'��t���t���}$�#ʒ�1�fRT�6ou8T���Iv�j⚼��Glp���TAE�k���s	��+�VnXK
���$��`��H����	�_��%/%
��"���J�x����6C$q�4�T yE��r�3b��������^��Fб�p�Z�?���������#��ѳ�ӿ�X�a�牍�JoQ���G2p�o %J[W�,eo�:���}��CMJ|��`7NTb�7>�jO�s�s�B�QXҲf�!�=��#V�V�\/���*阃fvӳ�
���G)&��c�@�96��S���A��*�X�t�C���#�a�13��9�\�k�?f��M��.��L0��8x6u��W<܅~��{�<3��LϠ�6�=�v�[Y��Mw����ki�N�`�+�G!q���4��(r�@AmsV����)4���ǵU�d�w���:�04���M�/�#�f�֜@�w��b���O�Xk��
K΍�-��N�R	���VX!�>�z�ԫ,,�C�X?6�܇�ra0?�UP�uN�#e�bq���>�$��پ�~��V�J�<3׿� ���"=���A��1�G���5o"G��l!���q���ͨ<U��*o�v]����d�l�Q*,o�h�\*Yd��b�	�m��:�?���MԦ��1�M-�_��I2۔�����Pl~)�v��5f+!!Er��h�+z���|��7�ن����&�`s_A )I��{����r�Vޤ�JU�L%���$�����A���K����6bOd���e-F����0��
�m�l	"Sk���zo�g�7�q��N��Ĭ��V��x,����F����+j]�ڭ����9f����p�;�U(��hL�<�-�Ȇ��]K�Kk+lJ%�2��*�@�N!}� ݭӰ#��Y����i^���Ⱦ�8���� dy"���U �m�(X����{��n�z胞��re�.V؅݅��5�PtЄcax����҅��	o̕�p�����?_�ߎ�9��0ȇn���� si��z3���7Lo��F�Fͥ0;�,Ѩh.� ��~�e��`�Um�~���7�Q�:m�5�i�8HFI+I���u��=/&ٴ1�1'�d�nCmFֲ��T����7�8��xǡ�x	})�<b-����&8
"jV�1G��.(v0��u�o7��l����Mp��q���z��ﾨb@UE�W��m5 ��D�|� �k�C�c�"�i<)���3�Й9��Rw�s o*���[��xp�ջ�@�#fs�S_d(Gm6���pp�P����!��[�^�=8��<-:l����,�y+�j�"�.T�����G����F�v�&�&��\�,�|���>Ch���#����R�}J�05k��B׬�IE�	��PD�$7}�_�ai�G���0Tr�� 8}ᨈt6�O��!L:�I[-���Y�bo6��Z�z�b���ݩg��d�l��5l����ʸ���Ã�4�!,'�Кo	1�m@SQ����C���Ŀ|(�����I�`v��X�JgYŻU����%���mF��d�|�ƪ2HL���W�<��S��_t"րs��E�[�#�hOw���c�GvD�u%�rB����g�R�X?[#.�Y\~b\��66�*k�q�ܞ�3)��m��(��k��!ݝӥ�/�w���,ռ�>�F�?���0a����X*���������\�4�V�}�6A�x
�h�:0-���`v
��pS����*xC�Q$�Ik�#+S�ެ���.h�]uﯿ`��Jw���m�̼�YyD3���:R���A�\�,��P��(��$<K'�KS��v�Qg�x�$�ڕ��b�;j��� ����<<�]��5�A]��B�v�D��ɫ\�XȚ�i�D	-�qủ�a��IPB�%�&hKc�5�7	d�+�e���	p���R�ż�T��PIk���?&]je���夎�R�?��F��m�}�^�ia �o�R43Վ7�g'�eK3s["+�JL[��	,���E���u��p��1(�����k���o�r����$-1�[��a����#��ەESy�n�/1]����V?7��a.��FT�z�i�)>gSD�}�M�W߲0w������M�6(�Fͻ�"�yU:���5��T-��`P�UXv�+}�E�d�Sub��wQ^�2�X��;<\ӫ�I�͗���<��6�B��R뇝m{f0�HY�k&��� ���H+�q��:=z�04UNN`5t(�e�ɲ�b8nz3�81$����JL���c;�A��V�[�ET�j�4�gnޏ��p�B���4Fa)�)� ���/^��AJz���ZvA&ނ��;!�rK���bd� ovr���.R�TZ�>N��V�`��WA�jJ
,"�f��Ҏ8T�!����f6o�W��t{�Ǉ��5�,����;��xW��K�rF7�\d8�ԄK_�c����#���M7S`q+�.Y����[�Ej4�
�BLR+BD<��-�.p
�GW��rR�D�ؖ�=��=�~��J���SW!�����-u�"0����Ւ�*��i	(LC|�\ݗIɓ��@��.�7�W�>-@�	�e�]j9s%�de9�M�`���>�_���3VW ��ɒz��B��k��)d����g~+ve��BBQ�O����������U��7x-d}=K@�Lt�n�K }1��({�;aej�d��A�|������잘��Sl�f '���+�N'�D�5f���Ac��j͹�؋��M1�1��l3h��Q�G�7cwr�X���LN
��uL���s�Q�3���p��}�.+���`�	i,��_2LO��3��"Z���T���H�옆���^����n0d��"��x _�yz=������	E�m�?`8Iu,�i��#gԙ�af/p��)�xۗ}���ﱧi!����*HW�E)Y}��-�oX�[��B���h7�T˸ӛ�pTD�Pl;U��U��������5ǯc�o� VEW�G�H+���Sv��|�/٥hIh�%����K��&�_�r������;e��T�;n��Ƹ��=~��D��8��R�3HYM�S�&�7��n���|,���+0����a�e�f�sX؅������֥9����3�O�����\���6�&���#���(xLH�o�\��{���>w��߸ܜ6l�Hon�V�տ�T���[�xI���ZYL��mQV��@�m_a����7 �fڪ{wZ*�G3~f����o�}*S���ŒF��p9�C���B��l�2���Ă�Ϙ��,>"��P>����4)K��ͬ5�B��q��_�+��h��oR �/DLME�jy��!�왌��B�X{P��h,n!A`���b+Q������P[TJ�����{�xdqh�ּO��O�����w[uC��b��P� ���B�*����sQG5S�5 �?oeNk�?�x^��/e��y[�s���1;e,���&�}0%��c8I�Zz�{l�7���V�$�ekD�u�@vu�ΥՈ����L�����������7#H���R)?�5^]6]mo����P.L�\խ�g�������E�']g?�®���	����w����K�6�f�+3���C)	�]_���}"n&��nͰc�>����!O�����_kvWA�\�4������́Q⚷�Z�H�]�r�l**���]r�f�x�R#BF�W�rJ�dʞB18�]57�pz��KK:�s�1/�]�u�Pg�pe�>��J�4ž�;��t�Zט TԨ��@|��I�^���C�>��WqB�9�>�e��j�$��Ҫ:;�"�����Y�����r�������[Y�1y�ť$��y=-�p�3*s��P����wm�V���c��2R����x��HR�̍[�)�z����
ǂ���@�K�gY��/�Q�����ñ�b�k�D5^����ɇ��u�%�/��I�FrO�6�/�Ds2Zf��C^��I�1R����$��	D��7wq+FM�3��SQFv�D�%I�m3�����6u�n�95�<R�߅(ip�ao2O�
�en������i$5�K���F�v��w`��v�����T˖	�u�^����|R���)�׳����5%���Y��!d��e5�A�CQ�`TPQzu�q��#�Zo*䀶��8~����b�/Iu�F��l�[�~�Y��>��k����G�4�!�_q�ٔH�cF����l�A�7�t�?��O����M�a��r��$�@��ױ��H|��%�Y��29=K�;�"w��+�K�x{��]��!�g�����F0.�>����]�m��O\2��>v�v&~]Z`��d��ᎁ�紷��D�)0E|�3tӷ+�:��'S��F�V����p5>�e@����U�WJ��]ᮘ?`-�8�ۗj�W�%ߣ0_� ��n�-�c˖��k]�*��n�D5���p��m�Td�7�i�~\�W��	3H(g1�R���r�R�t�8|�1i��v��h��r��W�~�7{��,��8��J���#�,��!Y�x�W��?�E��=İþ��yqf�7'��O��&<G�ΒHy��*�΢�7�{���ŨQ>,1Եg]#&��7��9(リ���X	�y��ę�̈0�jVJyk�t��<�0~�X��#�N�[�F����k3�T�T;�m��4Z��.�aP>(R!�U-O@D��=)�%^Ϝ� Ӝ�\gÏG�E؉}G�Aco�<���po�Ϻ{��ơb�y���t,��Α]57&|#�hj0pv<W6�P� ����$(�~�R�,T���� ���bW�2�GE���'I�`��`�QV�`��x���������3;^���T91�ɕ��̤r}q�M�K� ���ړUGc�D��5����k�d�㺵����z������ŽL�C�0Aj6�o�&��u�+�x���ȩ�V���ň�/��J�uS
>7<f�h�:.һ�e���J-�I�����d�zPi��ݩـN����Kn|S1"Zs��n{ƿ�-�>~���w��o��X��-r^�tZ{�a�>�{e&�(;7wl}ϣ��)T�]r���D���9��F�D�[e�}%a��؜�" g���pD�]�𰋔t������'[�/�	{Ա+	�A����U�A�
Y�Ο��$ŝH|VuF[`����Gu�w7]���zA��2E�8aM���Y��#������w�%~a0 A�Mj�gg6h�{45��O%��-��������	]yzs|ַM��If]�xIH!��+�����
��f�qD$��N���|Ǎ*p��D4�\s��5���}T�d*�	p�{��"��S���˒���̴�
6�W���p�g���
��?!v�E4VIt��o���=���[*���
+�lE���������6*C�h6
�a[�O�ss9����j�_N�.�9C�a��
%J�S�{[|�#x+��lI�-�$��fHN ���g�"gs�����,_n�}]z�{f,���9>Q.t
[P��5�m��O�7@��弉�˻�r�]+Q1
�v_ƣ�
w�b��TF�X{ʧ���:�.Y$dK�P�&/�N�a�.�}�<[]��q�Bvf[5|������	Y�jؕ^#o"��i����Q.������?2�o�>��־�J8�r��F0��U��p}эdm+�bL�s ���.�R՚�G��bM/��^������&��4��UJ=Ǒ�����4[;�}F����H夹i`�'�Z�o��5�v #M�A���|=��� ��P��H2I���hwKD��.e]���s��m��O}���o����3���9ќ�����4�s��o#�����X�
	m�i"���UP�.	懟=HI4ڭABn���r�����@㝿Gf��V�n��5��s���/�tC)G�R�S͡9�MWQ�h�T�	۰l� ��f���	��(����5�{s��&!v%�F��d�c�b�A����4�O��6�q�R�����캒�������M�m|�*n��C2Z��@�c_ge3�S��@���-�3�~6��i�]"2�Hᓚ�o�Q��@N�EGӴ�����W
��Qڼ�K�%�05+}�	���|�,�*���x����{:��(ei��A��o�g�t:��n6/YO�UJ*岗�oU��"�G�f���m��QGer,.������j�r_�W�IX�W��¿�ƾ�H�a^�g�yiH��Qiu;�x�.n&��}"�,�ı0�Շ�!V���U��0d{a�p���4�@����<	歋cK�����sҘ�d��%|C�>�~�5T;������J�W�Y���^��Q�24��	�^�SR�bS@�_Q�~ݛ	���a����˳	��.+?��ʛ9ogΦ.���젾7��e���Վ[�������j�#("����� ,U����gUͶ�
Q����H>�h�p�-+�RJaS��v�g�����2Hq��(�g@|��U�rk�s!^k$%�����;�F��PW��3n�W
b�*�9\��y�p��ݗݢd���|S�� t&��0K�	� *ٞ<P[!���h���𮃊���l6�|���(���x��>?��+�ǘ�Cd�-���6�����_P���}��v!lY�W{ ���C����Y���� �§M�Z&/� z����6��C��g%�`�a���o,˔~=�<hD-`�����h��XE}�8�kEID�x�}}�`���F�\^"�c�4���
�J��%��Q���Q��o_�	��=��X�� b�wT��(�U��u���EH��R�QbF��x�Y�.:=�[�T�����8|D���p7��#v5���B
�W�	�M���vz��6�X4�0�K��͓X�Z��`���B8�x��]]%gA]��-#��a���p^΁�W��2�D��O�k_� ?�����\[˧6.��Uy,W����֚�h�`jq�@%".
��'������h1�$ڐ7#b�Jw�����١gCb:���MLoy��$����n���a�o&��Ʀ���7��ډ3�X�i�' i5B�"����]��O[u2^���W��B�==�Xv�՟�Ȏc^���pqn�6�loI��&?�w��.Z>�4-[��G��|��W�+a�i���C�#��}└}�=Fku�Cm��Y��6��t�ϐU?6��i|.�Ng��ŞF�Oh���x#�T;��(}/���l~�O�x��g2#ş�>f���'��2!�D����%3�\���VyrhNd"%�'���2�Iw���O.����DYb�o�L�?�/JNl	Nn.�U-�hԎđ-�o�bh/2���z{��̀�Z9C����MM�)ly����McΛ���#N�	{���^�I'�c�X�{d��<���AY�b{�i��}�f$��b�,g��->�b0�S���i���LBP|Ș���P�#g�Q_`)]��'>��R̝����RY����8�Js�CI�����@M*����1��!�2~���க�be����.�j��<ƒ����3S�I|������5[�.�Hr�.T^P�����ټ��~�ߐLG ��*��a�X��ߓ�:�CNye�Q�<p��_� <�}�~��zw8�z51Ah��ߩ���q�vH�2�d����r��9:ߚ��e��h��+O�t9��n�,�Gd]�&�lq��D���� �AՕ�[���<Yw�>�L��ػ����v_�JDH�5�-�3l(@���F�4c���k��)�����,*@\�m�*"}�'boH?�Qc������{\o���J�'d���ѽ��>��QX�5&Q(a!���&�? f�����x�[��%K���N󲳲C/�e�a�˫eAh��VcvRn��oà�r`���ט��f)�i`�!)��!@K�
NHp�V}&��q��� ���E$����vq�Ye�i�2T#�H�J���O��\���tr�Ϥ!)��I�b�C9l��N5��
�����~����I�����{'����'�cD��P^N����1O�����ǋ��h������>�l�|�+�A��:bp���zi�}�̂��$Z���!��``���x�\{'C9�1<�e��KBL�̦Y�-/��v�Z����(��yx�5VS��;3�b���'J�D�w�l(�	����	*�f�= �cT��
��z��31.E�,�����R���w��n.G��ҋ�n�K��q9܌����^l`�J�&�.�iG�?x
�h�x'Kc���*6���<�z��q�#�qf&n���	��F�Ee��X4�>���x������(]���S���T�#g[=\u}})`�ko�`���>\�c?�k*Ѣ[ڧ�;��7��BR�Y�O+C�b*��>,w�ó�n]va]E���2ٹY�;_�w�S�YJ�^����4��'��.&�>����=�%�vTCi�v�G.)�XS���Тk[���[��
�"���vyV�޴���X]��@��B�R+^�L	#1{��>���JH$����������'��rx�����_ =n��#��J���_T����>QCP9��	i�+m.F,�d��]���w��@83�"��:bv^���DbX�-��D_��6\�?֒O��{�-^������f\I�ʞ1CX5m�:��	�Z��L7�Zl�n�FF"�3�<��;�*	]����a��Ru@W O���D�#A�_�7ε��T�?w��[�j�,�ѤNjd��5���A.:����mV�ϴ�v��u���G'���Q���n.�FF�_�@�X��1�&�i��=���\r�)���جb�E̬}E3q�_�#˅L���4���o�,�p����o�M��6f�a�����KO��nG�N1�Gu�
ޤѴ���"6tuJ�0�Ϗ�43�|Bh�j���[e�'XF�T�k7#O�)����I|Y_��}͉|��bE��
���1�R^����T0�2�l���sq��/�U@m�N�w���ڼ8�I��yv"�'R�EQӆ�X���Z�����b�2z�]��-��Iia�צ�[���we��i&b3}mKSb��K����;�8F�lu�E���$Vi����������ꓭ�0� M��qy!�8�Ӥ1g�V�<o��t����#|eYͥ!M<�hl�M�Ko֢�M��e�"�*��{恔�c�VGN�b^��H�$�=�ܓ.�m�B�@�}ü�`�/���c��3�]'��3�_��1�u��4���f�"j��J��<a:VWK��3���b>~Q<S�B�Ѧ�[s�UC���;􁤴e�Jp{�c�0��vO���1/����/��!C���d$;6�o�Y0$!���zB���˭��>�X�@��l�\���-�D����7��wNޤ����̵0L0�n6��T�>�	#g;o�Fց��B�-���o '��+��Up�	�ӏ����� e�GIA�S�(���p�3
x�(vf����C:,��p7JɅ��4�x�����i��Am3�zd܁���-K�Z%�aܧ�����M�Up�:�u�e���$:4�L<�(�ˤ��̭_�~;n�/�Ɗ��%�a����s�p���"��t~���0����;f֫mw��}�K��G�׃���Ι��8�{���g�%p�~��,��������T��?`���y�4P]���l@ЈS*�~�o�#��\��sܟ���|+�˧��ߜ\	�m'�lw���F��O7\��IS�ğ��O��;�~iV�=��OW=�t���E�1k��}���-�<JP��l	�S��6) �rb���3�vri��ҿJ���LK�
d�YWqQi_$��*���y��N_I����կc	��E:���Q���/)��Z=n�y�W�?���k��:���^�?�˧���ZI�I�ZyTI|q�.v�D�jG(�$m�]�_tR�`*��&�V�G: �d2|����V�KL�����PM3��-/�vJOT.�'uP�|ҙj`=��M�_���u�>cU���P\F��H,c�b�=�k���C{VK���R�14 [�7݌�ޟ�(l��aץQ��da�	�&AW����V�=�m�s�Vh���I�u|��7����)l����ƿW�x� �v:�)���4���b�鶿���9K9�S��r����r\�\Ĝ��������x1~]�re�u�$'r�w9,p�N�����@{�<S��G�l���)�4����Aɒ<�bG����H�ׅ�������i�O�/WP0�����s��%)�J�[���#�'�t���%���������ȳ��3I֯���Z�B�3�߉T�����ў��(-}��y3q��v�R��hq���K�,�p��h�5|�W���n�f����E�����LF��bI t�Y����s�n1��L޽R�޸$�M���A�Ք%�1ׯn�R-~�..��&���U���?��|��m��9 �Q�`����\��M��X,T�i����l0�Ŀ&�m���V���;�ED�T�aU]Kꆯ�C|������6%���ӧmӨbdpP�y �J���{�� ��?��~�]�`P�*P��S�ka�%��\�$�C3b�
���#.���fA��/�~ϼ�ZU^~��AQ5n���E�6�5>� ��I;�M���Z���x���B�prP	{�����IP��PB�3�{������d���!��Q�,�.<����^3�=��|���a�zΪ4�����2;DysVO(��ޜ8��g�S�X��Ы��c_��p��vӷg��0T	���ړq V��`~�< Q\"�+�Jc5�9ᬖ؆�aФ^�yi3`~"���B�qpUᕒ��Ь�Hy���]>���l��;l��NU_؈Wۮ�
��3k�S�q��4I��̅+�0�&Dozr��[��8��`1�Z�C`\kqt�-{ki��3��<o�^j�٪��=IK ��zL�,{�+ �^d&�}�lϲ�`3g.y�x���������Aar�Ɋ2n���ߙ��*Sp��V�-���{@/����m�ݝ�!S�E�(%�.�.��.A�l�Ǧ
������,s�"{��=���f�{0z��K#FKX?��w���7��NZ��냀��ӝ}0��^�S��u��Aㅔ=L�j�Ct��	�.m/K墵��p���D~"h���Je^*I,ֵ	�y�7���[�az
�Тb��b1T1s�۳o{Y���z���O㊜&��ѹ�6�61�P�c������^+�IU����ـr�W�~�Md�h�x�	(��^X�w��!�uz0#��]���>�H���O�?��T�j���l��okp�*�7s�LXsiK�l�-�������ǫ�[�bdc��!f���}T%�X�\�2 �#�Ts������>�i�Ѹc�~+��D�����l�s�@x��������H��u�.��]��d�sT�@�_n�3�<� �&,$_��b$���)�eU��TI�Uة�+�'�Y+t�+���h��˜��V�m�O*t��P^&V�{�Pk\�oψ?r��~�>�u���xON�v6-pg�j��A��j�{so���,d[���}�.���U�Z�������x��p�W'ʀVy�f�X�MBD�,�c���z;.K���~�jÜ=�H��-bUg���nd����5/���a TO�g��:��d*XЌ��	|���}e��Z�n�7�2�d
q�ٕPz�>gѵ�i�K�Q�G\�i�?�E�fgw�����mU��N
`�9i���8;�6�d�L�X[�)��du�xs��.���6�|�ሇ�|8��D%a��uݑ����*sqn@�c�ͅ�Bχ�xq���Nm�B�����\*�l�*�*unFl{�'�~.�u�J|�ĭ��M>@�\�3�	�D5e���×���@��#&b+��JXȪ*'(�ODïw���5g�|]G�Hm�sդ��OM�>��^�ʀ��m�AqJx�<���a���/��iQ�� &S��z��R�˪�
#o�IX�Z�G�x��"�#�M�����HqM��ʒ^�_��� �kвX����oy_���3V�#�A󹐱�DO���5.di1���F��[2ݭ�p�;�+�V\�	��j��曆4��p%�~��|���.tFH�����\������ʕN��'��i�^��c���]��䷭i6��YZ��cCÊK�>��� ���|_�t��I��?`��O>#PU���ǿ�6��6��-�	��n��dG/*�Wj��M���������N4	2�[UqȈ$��A�n�y�ر����!Ї�]�:��H�^�ѓ�{��\y5vlc��ڿo�^:0\�LB�̅(\�ߟ�:s�ֲ�_=�`d�w�O+
�܏��q��NK�8M�M�7U�+:|�q�RZ5��V���T�h����� Q���Hf�W ��3��1[��"�������
%B8����6�r�>N�#��9${ɐ����w)�&��[�Aַ�ԟZ-ޗ��ΐ�VF�l�sFW�i*5ת�f��sͿ}���ۜ^�v�d�b���)���C?)˵�֗���j�d�C��~�Z�*�mu�.��CEp���o�&�Cp���E�ӯ~]cE3�|��s��I���&7-�1%�j�{������:~�h�h�.�W�1�%����\&V���ZKa��	L�	��� ��?��{�
N�#�,bFm���~֔
���1�՜��_v~�,+�aُ$��&�iQ�T���6;�&�������_u��ǂAd7�� >�"
�'�i�k�US?x�k6HP�,����;�����8�[��Ɠ�_��rM����D�Wm[��p6APE0e�^��?~-�^��.�Z����Q�v`ŵ�<��N:��9�ي�s��s����cW����v�����9	�}BW�f����c�)Τ7��H�T\"����$ 9�#��Џ�X�t��{�n��Fn�|�ZSK��oP�c��|���rg��hJ���@~��]{B�9"FN��Þh�D���.s��x���ɻ.�����X̳�>ָD��Y��, _"����ElF��Q瀶�|`�S�#�u��m�m�?Q���$8�.�Ymτ��0L;o��-�:_��Pjw���c2�liC/����}mt���DG�o��S:QDVFP��&W].F�_���d��qh؈3���\�D�7�i-�!��tF]Hb�kI�.�8�&)J�®�I��B��0�a�8�@7�T�Sl	����cE�"�Z���5�v@=�V��6B`執44�Bz�u�V���0P�陣P���$̠A������l���O��L��n9֏pӫ����>9m��������ڍ�݂<��#�0t��R�=���,�aj"��`���xʃ=�(�M')�7{-� �^%�z$wh9�?��0*$�D�<2�9*��g�b�y�j����6W$ې�n��|�RA��� ���g�򷛻B6,����OLƸ`|�]m��0��y�9��؄s&i���u�M��¶ô���$0Z��U��s�ʠ<"~��#\>��e�7ƀ�?�a�I��:Rб�~��}m��	�e�W�Jq�KU!�o���M�Ih����*�!%���+�]J2�Xq��H���-Ó:�x/iu�H�)��%�jb�YW�)�D	\��<	��D*Q�O�'F�	��B�w��u.Γ�F����F_�jV�Yc�C=�L�oؑ���uT���"$W+^:f�qЯX^#������j]�P�ݬ#���W.E���.�!��y��28��K}��do��@^���K�8�7C�����?{MnO+i����V?����*��M�@Zu�#��΂�������4�Mw,�dK/x��;m��i�������#���ID
� ar{	�5`OY�,���z����AP�
^�Ζ��i��޵���^�W�<ZD?��,��p |�ۙ6q:͚.?���e����Λbۋ��&���l-��$^�`Q�,Dg~�PT#9���|���,�	ho30������!n���a|N���a�io����|���I��� ,.�Z�V�m\��i�|�V�k�n.��G��� �����	>+�?��7/?��;@��q��~�����4�b�cxv�Si����:���P��
q!5%)Vߜ�F�S�D�����1�.Z�nWS�=p���~|h,7�b.i����41�ʴ��@�jIo[MDb(Y�{��dT���J
늏3Q�CA���A��2�וX��[ƽL�(h����.�m��^K�!�%�UP{�6-�/0�!�~J��$�Lȗ��a�[F��p�c������@��8���e��]s~����(�!� ���nx�����̦#T��(�d�n=],'me*A��!g#�۷ޜ�}˟�/���,Y��I�Еq7��oE�Gv)���X���	f$�#Ƕ�z�����}no�K�1�suǎ~��4o��r���?������-�ëS���TJ� ��aia��&#女�?т���_<��?�y�[��;
������G��j������_�1�嬖fB��Y���<�̰7�Zq��uH�)u�c��P+5cIwYRݔ���4��r��u�ع� ��ȟ%[��s��c�/��c ��1�
ߵ��G�f��,2S]!���@�,�7�r��Hw��l��+��з�>bY�b����{�z_�l�!Q!���cG�7>�����E}�Xm���U�rW���![C��k��x���jw��%�����sm��P8��,��	ށ�λ7f�k뷝�7 h��ȳN3�ȥC'ºd�(���Ɣ&���:���V�e��T�(^�O[MM���w�b��e�a�v��w"�
���ם�9p�x����.���
�/r?k�.���;Y����)����
[�`Os���7kArzt�hfR�5D�UQ5ä�@��5���9�;s��M���ѓ�S��to�����藈�rAq5�`�Z��<������z�ʔ��?.��jnpD�+[Uj�H¾z@���*��� �-:�k~�����r����ѹ�}�0�ev@�=7�0+����OX];����
�6�S1tZ�����֊���Pp��;s�Rm����3�6�I��3wЍ?���cp�Ǝ������/���*t0f���%Pؿ������	��#�引[⧑ό�|0��2�&צ�3B���X|ć�J��0�~����&l�Qa�DN�t��K vi����PgQ����߫�s���ڛ ȗ��
X�B6�a([�ߐ���?�z=�v�'�~٥��BV6*oT1�V�/����Y��l�r�ދ�,dc���ߏ=
,�.�`P��@\itt:R%��)fm*N�`bĨ?~������
�#T�s���F�柳�;,ۈ�)d]<X�﷢��g>Ú���B�_�}��! ��͖����\U������x5�O� �x���P+�d�tl���v��4����I�?�%�W!��(oTAX�.�Wf������24�\�$:#�5����lM��qw��2�I�W޺��'��z�5����-�e��	m��_��q<�*���jIؙ��:�RT�Ζ���YT�t/�1K1�7����
���-��������&�DU��\_�|/���^0#T�����k�C�[�%�k�j�7vc^�LV</��} �W�k��:�'��D$[S��˻��HOlǴ���3���T^wR��IA��"�%fS>���"����hW���Cs���>)����m����p��D�s�])����'�y2���cfE�� ����mSh>V����"[I��]FPG�ݗ���3���5(�n<]I򱓍�/�Nl��v(H/f1�"X�ec��Q��iw���|�}�_�o��t �f�3r�׭�*��N�}��>�ƙShkȶT�I��6�ͬ�����Vm�������J͂�;7���]���1��x,�B���Y�*Qd�G"�;I�	���3t�\ﭺAQ�)����q�^*�Fj+�5[؃g�&g����CT���Gk�q�~��P��5*��[�����#]�E%-2J2��z�'�����xۙ�I`��݀e� ���������W}���;�r 5$��u�m{�Vw��ZX�*1�ʹ�cZ�t,��Mn~k�A����q�����ؙT!�N��2���������w�US)N�ǩ��2&�r�8V.h���/��Ơ���*���b #�ˆ@#��
b�Z~=��*5��1z6��F-p\�G�y�鋑���̝��,Uī`�'B0��$�`C!Z-�� !�'@����h�m�,D8�r���
�&���v)g�> ޗ�.4��QͿ��}{�	�I'"N������eE�r	qv����xC X����2�.�q]�l����/'[�vA�Z;�����)��B���"F8 ��h��.�Եe)�]�i	����֮� 75CW�,e�5�*�_H�3:?��{��9��g
k��b�U�m��.~�h��-�x�����B�U���+:���A���hώ���	���L���>$od8ؼ�a ��������ej�]��UD�{k��HH�ԥ�%`�vhZ3o%����9�Ł,��e#w}����<��ƫ�a�o�����8ea����}a�͡��6~��٣5Z���XnIK��l�v��}�ݷP�w�o!S?�}bO�x{K"�gMm���C���""*��.���b�A��d��$��0'fSy�xU�d�5�
.Iض�Ӎ��KYgBX+@��Zc�N�F���<����kV�͝ Z8�"&��C�FѪY��C�`]�ֹ�-���M]kV@ܷN3�!$�]����R�R��R�Hô}��H�O~��R	��I���w�ǹĮw3�@��2���р�ق<C{�VEԩ -���I��d;��C�z���9��7�ZJ����@�{���4g�A�!�±Ҩ����ә1���џ1�d��w��Uw6��*��U۪鿢 )1&)�Aj}%�q����fl������.�����HOY M_a��yvΘ�.���wϳ�����}R�a�%T茊_![�<A�\��C�����0O����b}#j+���Qjs${Hk{�A�ah`t�����-J�TA�]&L$��qء�<6�N�'�D��>A��6 &��i�((�pU����KeF�	Q[�8n=���*`> :�VSw�F��H{C�/Im�����ʳ���o:�����E��h�{�9�.��#����-���g���6oФL(U]��q�U����W����RO.�6:9¼���ݎٓ���N;���iv�T�,�.w)��u��e[��!���d�/1_Q�oYg�2��lB��T�Ҍ+�>e�n�������c�~i���Aw� ���|m�Y����#E�a~I�T�X��H�:����&W�?���_~]8�xT��88ќ:�'�>W��H�绩�C&�x���K��"����Gܽ8�֝��J��f�\��G�F�,�`#��,3���"}���r �2�@3\)�vxf����]I m�$IN"M�L=���8�"�L��}~��e|������ם��-���=2�_��nl<���'�)���p=���}mB��\� v=K%�����G�}��U��E��%D�v��e� �W�1�/���f7�ύ�����̝�#�3�'��1�k���u�0����:WBWH��.^1a��C��K�Vk����d���)犰��췠��f<-w�~��8=�����x|'��T�#N�@  t���:pWa$����V� �r�e��tld��X�p���J苪��#gg���At���6��C�mN\�P���=c���=�4���4��q�����8t}�2H�<�b�w?�$��-���EDb�0�L_D��F��u5�BZ�:�\��a2/�����o(�]І�ɂ��cFE�{� �g�c��_cO�#��Y�0-F�`g����[I�V�g3�<��T��k^�t0����QJ����y��0e�&8ȩ�z$�80UóU��OC��b�'ԏ ���:��WN�|�y�0����~�b�D7XV` ��>LW(�����c���{nI9deu����[�%�qC�JYl��,m#c��"'�L���J!6���Y��[�4/読���~������m�� ����ָγ�8�Z����L��0�%�8E$�ϣ�K,B�P�ٟ(��b�{�m�l�:�;�_��ݓ��k�X)cx�Y�@���Z�,��W+�@���A��^v^GI�ݓ�w�ȼ��l/X�6���Ĥ� ]4�6��S|l��#���K�N�n�e�Y�Bs��s�5@��R�dZ%!R� 8V�r�n����x����$D���];���xBO����W)`�\J�1��JU9c�%�����t��VV#�����xE�	|A)n����Mİ�f��3b�,g�+��K���G��P��a�D���O��F���njڶ�	�g�ӹ��؎b�R�'����K'B�e�ʻIx�W���x�%jp���M���_�Z�Ξ��m�A�6�P	L�S����>&�Q>f}�|F��[����yt;Ă�=ȐP���=Vng�D#!s�,�m	N��^a�����oY�d�f`����K��S%U-�/,����S���!K�B.`ɚv��p'ΑC[R�?��M6���2G����k�Pu���!qN �����v��<��"����~j���ɓe���؅��sW�yM1�y�����p�[G��ecT���@䊘�8������=o���Jƪ����ܢ�1����G�>�W?~*-s�m*=cA�/ 4�8�H�7��.����F�'����/o�o���Yi�q����%�����E0Yw��TH�^�$��GE;��̈́:�?{4���\�m��^��c
M��E���t�,���nY�$i��[2Nu��JS/�q��+���v%����a����880h��wLG󠻂U���R����\�wꄫ�H��K��\�7�������a�Q�^� �*��qy�V:�< 	b���ﺜ#k���*��q�vd�wCa�#�
�%��<�r'ҾPYI,p2�o������V�ڃ9�@��\�h�7��ޗ����(��X��!
�OE7?�>
�&�s _	Zm�k���ڒL����isP�{���
3rxj�����D�R^����*(W���h}/F���r��?��r����o�c��w0�W�K4V.m'���r��̘���Z.�l�g�e�X�Ʒ�����2����9��Z�d�h���z�W�:K��P�*�@g���'�G$Z���-`4�cE��;͔fh�+}4����+웭�Z�/�|�'�(訡�(�8m5d�
�'����U���؋%�H��:�K��A�J�κw�>;X䎖��kk��4�*XAXO� :x玴��Мz(�ӵ��W�:�%2&G"D.\S�#G@�O���,!,}���e�j����� ��h6�6�{��d��!�@ȴYL�+ݡ�ϵ/�r{Y�W��:�3�q5��I����n�QJ�MR3j�"��?�-I��]Ç�E0
b��0�8�tC�������������c3���mw�(�8���ͧ��/���jY�{�v�)Yq7Jw�c�H�H�Y�h�i��F6��s��	&����񔼺r^WS�� wni��?���G��l�[L�!uiAi9-8;�M�gsB��l�5�
ر����&��'�-|�~8��#M�`�S4�H�}��{rv��}��n%N��RO�Z����Z��槥�S�c�h�<�;L�	��R~Lhm�X�ǰ��T��ZNǛa����ՠb�.���~�(��dؤȈ^�f݁��VJ�_α=H�LL�c�w ��L/��hq"����cqn&�qc�"�'�V�7��4�\��$̽cŚ�%(|�+�!��jB���I��Z�]Z,i��}H�*��<*�h>a� =~��$bI����/B%�"p[���S�g��]��I�����~�^�」t�A��{���]�]$��/	�Қ%k�����s�����Z0�x��C�Dt�ȍl.R&������=�3��u�����f�|��[װW��{1��16	0aa�[�<� MBm���܎�*M@�H*!��c_!�^�[=,����m��Ŋ/mz�n�S �?
n����o��"Gk�_J��H/�<GiE[~�~{V���E�E��E�6^
NE�[<���B��<�i�#�8�!v]�i��=���D�Aa�hA[��`���YN!�(��ċu��H�%�b�@��=L�����0� ㉲��iB�giZ��7ًVK$N!���WXV���a~J�d`�L'ɭ��Z�5����р#>���UG�K�_��\�%+r�)�1�S6��U�{�S�	��J��X�9G_-y
��ʊ���pǂ�8�J�-�����){;�~� j}��*(����#�-�}s�3(��.�����������Y�|�2?2Wh-/��������%�z�-�M����$ݔm����Z��X���%R��J����S�EC��#�ˤ�"3�r���k�B�7�n�ŋv�$��͸���j\0�8�������_Y�q\��W�c�E�q�޿/A/�����X�}eZ�R�4ݡF��c�Ll��w���OBaB��X1皫sŝ��^*���"*�/:��[��r&D�ܭ�6N�)�C�-X�"���n}m�yO����s����Sa�D�����pc�35H׃��|*�Ȗ�(�y4����,�e��J1T'H2;���RK�U̇DG<��R!��+�N������Y5'͵��{�9Ǡc�ar��`����`�5�M[������E�'���m���H��D�)�`���kL���\�?��F����L"oӆ��핽YV��CV����q��<�B�9�_u�\9�A�����R�Țn�Y�─�(��]3Bj�P��T�>^wYM��d��|G�r�H�0�%�N���yi~��4��IG�}~�[�H�̘ ��/1'�a�=������Ju�W;+�e6�e�o�0Z�xoD���q�g�~����A�qR]~i�K̩�߲�3D��l�\�dz �<$���"5`[��ӆH�R0Ї�YG��@|-���T�w�?��,24�W�(�U�+���"F4︉�`݉�;��5��_ښ1��$��d�oZ��D?��,U��
���F��@���؂��<�`�Q�9��(�������K�m �T���ܓ��&O책��=������b�p,9?�� ���g�k�(����ctF�x�E���;��2���N46��Pj��Ѡ9?�����l��ٞ���0��D%۹3�L�o��F����Pv��T!b������i�W�,�M�8׻��	q�aP�"d+��̘uMz���f�hK���d�wl��AT��"��;��*�	�}<fm�{p@��^�bB&�` d��"Z�-j|7G�z�t84B�;�쉭��$�Й.�[̸(�SC!��]��'�̔��㇩|�B$�����KF��yBV�q|����;�c	?hF��u��9+n��q��&�1N��(��7��S�gq'%�`)͙!�W�l��A�����Cn~:K�u}���f���!��.D����NO���,�=t���q����S][-El�t��ˉҫ<.B�+�f��8��T��|�4�o��/"}���s�bCˤC��*��8�I����|[�~ߔ]P�%���ah�k��t$!�G��7��������z#x+����6�0�Ɉ聄Ч*�����1[
�Ix%&WQ��0s!3�K�Y��kY)�Y�C��FY���\���8}��[�Zf�]�_��Z�$Nz�֧\�|)RKg2�Jw\m��������m�A���z�e���G=��(�"�T
Fw?��?�	06_�R���������K�U�a�+�w��C\"g��63��>
��6^uݔx����_ՙ _�클�7>����2X݉��C��nc�[:8V��S��BC�EE�p,a��ł��=0n�����)L"�v���^Ħ�g��{h�h���Bi*��.�M �	�e��w>����,}���C�*(;���� io_���;P�k7ż�ք�6�,o����[�;ك��e���r{�}.�Uh*����k/�,��;��6y�:w̱{���Q����G�ĝ�<�n��ʘ�*V��XO�]���c��>��<�"��Fխ�� N�\�YJ{�Z`+����pΘ�O|s�bvW��P��T���W�Fz�` �Inۜ��Ӕv�9�3��I��w���� ��^kϗ��\�M���$P*�e��-lULd;{�'��PzV;�<T�MO%x`D-f"��F�&�9���"�������"�Q{@;��Gϡ������ߐ�r���@�6��w�ڡ���a��P���Vէ��e�٭�~e���9��ɥ�Y[6M��3��% pP������xC���$\��x�G��a���ݧ)�����HwBqE�|���`c62J�V���~����C�~�?�Ǯ���$T�:��z\�F�{4��c0
�����6e�R-�{����L%?m��Z߰Gd���|�w?�Br�/�S��j�s���
�Ȋ��� �Y��x�1/>ϺZ-����eI��%��oRl2��T:l6Ƌ��^�LB(k�S^����Z�@%kE�|<�l0��Y�N[܃��l��nxU\���5�L��[�Lg�mr����m�[+q���Q��Bݤ�.�VfH;��kH�����T�xrTQA��co]����1�����ܲ�e|dR4�:X˙�����f64F�}��\x'��\g��Rj�q��TH!���N�R�)#��=0���F��j����r�#�Ƃ�u̮Ƽ&#L��Nn߻�g(�q}(�7+^D!�׆ض9�_�cK�V��}cI�
�) npQAY"Wշ+�P�2�%���Q��ra=��e?ܗ9�<V-r+8j�S�([��
�V���Gs&ZϦ� ^� ���XsH��9;�@����S�D�z��z�m�Z]�!���B�����!����	�����)>;N��@--�Ǭϝ�T���ό��ݨ�+h��N8H]�{�����m*�ZSI���pԷv��ڞ��s���
hgt~b�/�_�����V[�-�1<�]�C�[�,�Rˆ �Z�Z�]���	�2yͲx��U�9;o��d%Sw]��mH�|�J�zH�e#"���ن�x%��ZjJ�U�����Ot��A�; ��������Ab ������J��@��(�����j����l�z/�]A?���::�5��{�+cH��=��]N��`�r��8�����y�j�ܘt�@{0H�ꝛf>��F�"�a�`���Ǒ��7S�!�G�kGH�h,��~��BC)��}XV�qnda �b���)����갤��:ʘ�$����7}�;Fd.NRN�H���/Ԑ�9�hmύ���Hw~UO�����;�VSA�t3J�,{b�A�����HF�� ����,(	�_+;�/ea/#��k��73�b�pƞKS�H�7:�)��ڳ��A�i�(�%� ��7�_��ņf&1�7 G��pܲ��X����>���O� 훓2�� ؈��L�nZo�n]�-ˋ�-��={���2JN=|�X��/6,���6/il�A$a,e]�-MQ<F��s1�pr�f���*9��� ���E&�8�.��ӯ��|�=$���T����"�*��c�H?���@X������ƻ/�V裔�����}J�QV�gR�ȁ��#��C�-|�Ω��6Sz�yB��������0]�h�2%[6t��e�~a������-�xic/�C�6X������~?��]n�!�@h<"uY&h�a� ���&e�?�k��1���LA�5���L�Б���Ԯ�F��,�.e�&�_yQ��蒪Ӊ�b�G���m��@߂4��A�ą��C��oPk���2S�py�7����\�8�jlV� r�ɮ���W��њmj�}�orC�8`i�:JB��I�f�	Vo*7�-��u�J����&��y�����!Ρf)i���{������3�_㣂m�p�y��˃���(d��Af|��AGu'�L�2��	�y>o��қ�ZYUϝ0/�?(���a��pko]�FL�Hb�b�2ΓX��Q�����qW�!�����e*$a3N���bzf�C��̸��g��Ɓ�5Fw����"	��	6��xX�j�� 7�<�p�����HqE!��b����!������>�ϡ3�2#�2:�Y�?9�bF��u�������^."��=}�s/+����A�$�4�w��O{�5����ί��!�}����5�e�H����*����	Y�j����OI�$�[�Ή�!�*���\���8�� r%���$�lV�U��Zo��pO�{���Ib����- �3���[�2o�,qqg��zcj�1Xz�0���D��ta�R+�v?�0�]Yy��w�ٝ
�`�J�����4��DЁ�upW:�My@^�8|�O�y65Z@V�3��ͪB-��������;`��޻��+㵡y�k��g�<�g>�CB�'�,�� ɾħ��O��C�N�iNo���۩�bi�a��3h	��+:�2c��>�J�.������O���b�\���C.?��{i�����d���=�O:E��jgfX�����v�!�:`�%�u~�[w����|WڭКzvސ�D/�"�vVb\�d�|4��d\��$VxG��G�V&#Ny\"��Y2	.�'@�	樋����j�i���3�YrN���{�:!�i[�'�rD���KM}'v�YIH5�~��R��bP�2L���T� kx4��PX�"�õK��%j�ͽl� �摱QsQ����*
]�.ɡui5�>��,%�W@�H��F{]�I*~����ss��¼V�kRge"���8�FP�4���Y4k�&����@O����n�y1�OnU������T|����ۭV5��]���������c�����mt� I�:0-U0p��7�eO��5u��'"ĕ�ߚ��kT}tEWK�A��M���*�%̬��OC,�;g1���v<B$�Cg��W����ǵ�nr�8�\��j�%���f��~�JB���@����GJD6�!��+c_)v_��eE��Ѧ�5k�N�U��뗽Q�NW���%i�S��Nm{Yz�J����L_�������0ޑϪ܀(�q��o��O�o<:pv(D�rGbK�Cu�M4q�D5'��ڃ۷��C��t]\�z��@Oz`�g�����c[��U#Sc�n+/��pMIk��J�������QCBEr�����K��@�"]%ny�_v�6���}��b������A����B{Ї�r�	���q���|����������F@�w�H�ɲ7%Yj���;��^���(9��Ӄ����^���J�8��J��;^�� ��.W3.o��_�������mދ��Al��G�[�8| � �E���r�	|�4}5?l��yW��ZR% �q��� Y�Y��x⚪z�@���5&���4�-�F~�8+YB��e����E��G��"����uJ������mm)�
^5��N�L>ie�}�,��ãb�Zi�*]�  �M��`����e�쭌K87$]����*�������{n�!D?d��+�	E3bo9mT��\�OJ�&w�*��B5���@|I�m$8�l�sjryDMD��&�Pۺ2m��&-wĀ��:�V%���zܰ�>%0��u�蛺G#����챋B���1(ө"�\�\X��vԓ}N��0�ֵ��V�Eb m��CźG�������?�������g������U	�0EԱ+������('�ڻ
�kX�� ���tLg�TŁ�n���ȟ<������@�V�� *)L3�7�A_�z���h�"�9����F�ӟ��M�ٜ�P�N
`�F��9z�+�#�I���N)u�[F�kF��S�,l��LĿ��9��r�=�z?c/Ux�^�`��'�C���E_!+á���j��#igIꣁ�������߲4��H#�TxΒj�ǚMn$����mn�1�%��K\��H-�_�_?���Oꖥ2z�u7�$LA�£g���H�xƆ�3�����8���]6����#��g�ݵt��8	���hj�Ef���[t��s��|`�(،�J�9��[�.���$����7�n�M̓���X��~Y�P���g2k2�)�^+%�wa��G�J��>��`u�"IA�P����zs�!m>B��)�:Bx�T��j8n8 �CX;}_�\u&\a�����i�
��XVKj��V���8��ޡUs�}r��C<�xA��l�'�[��;���ί�^�v���U�+����=
��v�-9e���,��̝��(���nYع�s�BF�t,��a^a��2_	�Sp�*�����ܟ|-�̠��'>S3σ���0���6?��S��W��+�?���A|jڠ�ehq�����Jظ8	���}IA0	�����8���I�k/�x�JjF��aa��گHH{n��mq�/�ܴ>�˃_/�ѭ�Y�GӉ �~�G��bT�ˈ��l�����l�Ǯ�yj%]��+3���_V����I�Pm)���T��56Q��S���:aq!E�oT����sh�?�ݖ+�Jl�`���8P�kR�cY�}�M�@Pl���'�"tA(t����\Ѡ1��z_���SF� ���w���j0��U�k E �l	*��cG�=X	b��/��%~�	�%P5���6���
�т��D�&��l��9�ܷ������ޒ�Nރ؍�;�s7�1��9��I�'���F�~�gl�#REr~'�-��8z[��l���<'v�S
��q�F�/m/�WZj�N���5gTǽ]E3�H|89�r������1b�I��������/�ܢ�<FL�5�4F����녳�7:�<mj����jdAO�����L��<O������v)��5C���,3�h��\���u���mj�]�n�$G�p��?�dU��;�5|�=�&��S�W&����V�8�:k������W5�P0 �nڹ=�4��E�C�X��#�ډR�s�%�9��5)�`��K�?����C{;0��'~��	_��ɝ�z��s�TS����Y+|6D��ճ�b�S�+�,�8�Q�X��"�k��c�$�}D�'�	6�X�o�ʸ���qr��nCa�&�	r	���W�4�
p��K-g���d�@Q�h�p�������\���\��҂/�R�c�����V&b��*!��k�a�+3�1��v��К������Ƞ#�3�ͬ�7��tf��>�T	L�����U�y�0
�*�aMQ��>��0=F��.)�ܐ��U�7�߷��@/�����<ە�����T#�U�{CJU\�{d!�gC��E��(���&qS]���T/
4#������v��cJ���só�0ꓨNG��s#:�J�Qv�1��n�z�|�xJ1�o�Oe:����D�P�h�h1�5	�SJ�W�_��)�|r0l���o1�&�M��8Kj3��Ab�31��z!��׳,;�aE��dm�����s�}�K�+���f,D��0V�.��"�ӈ^�������tt�n[%��L,2� ��<t�|O��}U~�7#@���Lö�i.�C��Ps7x�FAY����B��s����(>�G1#�e6�\�¤��Ï�>�_P�� �����)�����f,E���q%��S���o�}Fx�x�̍Ǌ5�e��ݻ� <�\�ږ���~���mi.΃ݍbm,�?�7�^O�誎��=4"�u�p��~���k����F��\���| ����¡9>��PP)��Fb�m: ��O*Z		��[sR�)3�zN���8*���<k��_�n���g#��Ͷ�����|ʪ]�̆���	���ѕ�+6�Sղ�^��,���t��F``������[��G�:u�4��ߙ�(�O��>X�T�HH�3�e����Βt
�1hY�ٹvC a^#*)�d�zD^S�}�*�����c�5�0�s��M�*�k�?G]aװhǣ��)'����gH6J�z%���U�s��� n|�L��0����)���d]���X����y�I𶞐VQ��7A	�T���/hSa,tT�}��o8�\���	$W��ĂWt��t ���p˥I}�W�I��K
�D'}������P���gL?�-s2d��uN��{C���`��*�q61t���o�#ekS�OhZ U �.��W%_�����G��㏟w�sON��U(�:�D���}�����dQ��������W�A�2Ȩ�-55M�Vvf]�GAY-Kؿs|?�{�5-��J�9}[�d�N�Bx/��4��=b��5��~qF���z�3t+��@�Mz���W��fn��IhRv�r���3�B4�Y'�}�2����QA���C�C0]��1 k֚�as}�\��xc�
��_W����l궗BdD&� ����ɏ�_(kG�Nt4A#����5�~̇�izc3�ŀ2u��Cֿ?���2������{޾��?���B(HmT�?���<��p*�1(�V�u#di�v���H��[�+m�ކ�4�w�a�7�_�q�^��9��9�͸ɩ>����x��ɣ�m#�@����,ȸن����R{ܭ^���}&\�l�4�g�I"_<665��!h�;�e�x-�[���3a㯚�������5Q$�Ts��p}D��"�H�i>�	��h���ā�6}N��#ՒoV�'�R|�z^�j��3:)xt��L�aJ�������5;l#_@enb�����h�����yq��Ӯr��O_�3˰]�m�I����K�T��zf��~���_�2V	���&�R<� "u�P��~�F�p8#í���4𕴗�`mKQ���$� ѿ?	�w��AU�V�@�1���-;|ֻ�8���9�x���T�.�w�+X�	�[���"�5�!�)����slr6�>_��7u�ۀ~���K���uTKi�e�R�{�Y<j��̅��Vܥ�6��Ch�/!��gd0;��1/��x����Ř�u	��lҾ%Yw:#�Ҥ�`��;��GmcX	*�򴆕䧤R���y��!@�|.�U
<d�!l!����+�ZB-��c�(�'$S+a�i������Î�,��4=@��p�x��}'���nD��%0�u3��'%Y#��|j�
�)���Ww���pÛ ����z-�;O�:�|�E�v.�T,����G���
�ni�Ge���Ώ%b���i�����su�}��Y,`<���ٗ��Ƃ�`�{���D�9f�\=��c��D�i��V��{����Q�He�݃��aa���?���􀵤�U�p��9W�A�8��$34ޕ��^����n��z@��ȱW��#\_$�5�dʰE&!��R����7�!ۀv��'��#V�y
Oj�ۨC�ņ�V�?&/�Y.i�&�A�Z"6�!��7z��v6���0�{�	�57�E�W�������l}���,�7��tP{k���hW�Xt�R�����ICt��F�5�8'��߮^���^&4Ļ�꒘�^6#ݗ�؉N��7��_�U2���]V��?)�C�ߝ����]_,�4�17���v����#N��~n��!i�0�J;�BO�J4�qNc�YQ�iM�7�z�\��B��K�P����z�'��Ȕ�k���I��$�_�p��>�B�T�ś4)�� @J۪�e��.��=ʟ�u�+7�+~��y"s����qIG�!����mK<B�u����Y���x��.��ݬ��W�u�o�����m�46^=.���"$B""��i�f�e��-���dJ:�x܋�{�u�y�v��+�����1��paw��)M$����`/�����nf�MN�"Z�ʌ4�h�x�X�E�U��N\1\j7>"���Ri�a��qV�(���()l�=���]~��Sҍ�n�,·�Ɏ��*�^j�D�s�1(��ʴ���,�'{�}J� .:Q��4#6��SAG�ȍK[,7L�����`����
0�by�|���p�p��xF���݇D��x�ɞ:3Rf��0C�)+�<�P�<\^�c>��*�U�ɧ��&�BH������!R�$������n����+~ĵC_�J�&�� �zf��-��嗜�J6|��u7��Y(�u�d��a�ۼ�� NpTB�,�ܨ�?͜�1:B��	���:���=�K�l��~	�C�{���7}��%�C̆C��iя���/�]���w܇j��E"�=����;�����͎wX�l���U8�F�>�g>D=uZl�*b�#��Ŕ�[��gjY:��,��B���m�>��|O.���t��95�=�ȸ:��vr�jҕs��P��jX��g��p�����W�;lX\�cs�l_j@�9���|VgAo��[Bj�V�<��������&y�8��E��Y���v2?��Ծp�@�V�~� c�G2��]��J��Ky�y*%| /smCf?<��kL��_A�O8x ݄gu��4�@*���a�m�����?�7��=�sc ��%��w8^� ��6i�tQ��N��r���qkfE/���"��u���g�m��ar\�!9¿9�qe"��WQ�s�fl������S�(\�м���F�8O�j4�7�JP�A���rD`E��bS̘�����7A���m���o|�$�fk��-xhr��Fr �U�����j���1��G �É�02+��e>���>�,�tu17A]4�_��AP-x������AܜWE2������+�̇@���[�s�c��4$��nW� �10-�0M�(�ѷ?���'[�ܸ��>��A/��e*s��l��*{D֬��rj�Τ��>�g���#̋��&[�� ,(]��i�a��B�b���1�F�I6����:kwQ���WT�h�U^�8w%�<�|x�Ÿf�V�Ͽd6��	qh�뢅�֒�t�D�ĬQ"^�h�u��Z36ߥ�,lX�)�M*S)�4�����Q���	���	����Js*�Q:ᵕ�)����s����_�9�B�US�F�is�jo�|�˥��	�O�[��B�+<��-N`�|Y&�;���R�.Sz��v%��|���� &�H�۰8d&PO��Z�Ţ���$���ʲ&�|�:H� В)���e�2��Z_���q�;����AY�U;�r��7I�[�"�{���˄���c�`S+�A���9=���F��|�v��ǁ7:��ߗ9� *9��^��b(}��硌	7h^W��H�e`�>E�W@�ޑD^��?���ζ�g�$UQ�l�O,��b��J7�PF���;j#����V��;*:�V���H��?k��2P�M2�c+!I������B��Fp�t�	Ƨ�i*]i���V`��t޲�L0\i���mO_�r���j.���g8��o�)쏛�H��9��C�w/�rF��Ռ�,'�wrEO�R��@w���u��[��I���.�*ܹ��$��_=e����}���p�Ɉ��O�
qy ��_�$_�9�DH�k?f�p�����7))��QN&��%+�>Ά��4��GDX:�q�Hr�s0u���۶��h�]o�ӏ�x%��%;F�(;�|a�D�q����cw�w�úΛ��U�Z �nr�,�Bpϥ�Ã��b=��p�W��Kz]
&��(�h�|��ו���N���c:{x}��Ptj��\��޼����mv���l�?`Z��m�)��mG����ڱ�W��Fg;K4��>�БKP�4��᷊�um=?��
����'�ɬ�l�U���?�G�K�w�N�y&��>Q�r�L-S�Z] 
i���ļ����������<L�\���w�Չ���Ȱ \4��.�g�0��� ���2��\x�2o��Ύ�O�rY/;u2��@����e�p��*��v����ʺ�b}�_W!��-� -&S}����0v���cg�h�C�Wm�
U���Y��}��	OL�x�o���q�9�{��4�MqT��[�o�\F�s~���E��n"	�5Q�����j��cf����
$�vw�u��������0'6���p�D�g �o��(�P�ⲻ^���t�@)���*&���{m8��G^j���������&���sU�V�y�w�����x�
�S.������=���l�*�����1�>�_�c�v�B��F{��>�m��&.��j��[ �f��>�����V�o�v��M��"x3&�IB��E�g�:{�U�e�@��g�ퟬv�����)��J�y
c�cߥUа~��){��t��+��mڨnr)�1�C��Z����9nΙE�ze��+�)8����=;z`]''�u|*����+��/��}��s�N���~���[�������.��$�}ًב\#�!���j���z�`냘\���o��% 3 L^So�~�xqKdV������qo�$}YU�fѰH��Wy�3��6�RQp�S�I=���b_�L`�E�o/ɞ���Z�ʠG �P���a��U�K�'��(��-�UGwtg�)��T[���}�1��}��lT?�V����{EZ|Ӊkb]�g��t[��;GZ��r�N��s��hK��[��Rs��N�Cy��(6ТFg��%�̦����}T�q�Gg]���j�(�t\�];}̘���Nm�����[�U����j~��ha����f~��Ȣ��@�� ��S�O��Ș��T��/TJz����.!�eN�y����|9U�4d%�܁I���a�n�����n��J}��D��Z�m����':��g����ow2)�pL���"�v>s�N6�j#L���BV�od �� �:���ql�-#MTd�?;5l35 ��>%�X�K"�y�,L(^u@w���aT�J?ssGmv��`������n�*C(j'~�
u	<���U���78���Ï.��yhW*��$� wձ}�5��i�镯=�ϙs��,�x7���
�.A�%�n ��v6'��q�Q��K>�Iٰ΀�������������~&���<m�:S�;T����!1I��Z@�4#uݝ�� ��W6z�vD��j��>q��p���kF���D��[c ����8����6���su�:��G��{��9���a
���}���!����á�`_e�Gh�����li��jSIc��G��K�(��Χ���9\��SO���|�1��=ݽ�O��~ �8 ���r���Qh�G�՟+#��"�����ґe/\�=*�����@'F�\�D��6�i�|8�2B A��nj	t�#�5�b��V� ��8ieO�ڿ�5;u>���_>�
xsKX�
��X6b�웴���+	F6�cN�B�Z��;��F���vx�;�	t猡L�
�^�Yd�Ԝ��'�ӁO�J9���L�-V9��2�^`�s�	2{���t(���&����w�y;��zK8n�H����i��4.���U=~B�u�4�o��n��W���J�}횉H�������Ͻ���{_U�B��GxcIbhh����l��!k ��67i�=H�WuA_�$a�7�~���/�r�Vbj������n�jN���Z`Q��w���*��F%�Ch��w�<5y�"D���p�`p�kP���$��е9rY�V��s�`a����"U[��h��ȓ�*�.���FT� �:)�}z��Teaj�7J�xw�r���ݔ9�̼�x��E�k��iG�b�o���
��̴ ��,�aw��9�����z�����nA�;��[0�����D������PE�;��f���.���\�+I'�Շ��p+��|�ka	�SYR� NQ'f;��'��s~
˖}Kћ�B�aA�-�x�9���e�U"}'e��'\��a���;S��>(�������&0�Aￋ���$��M(4�?�f��l�b����X��;�D�3 
�\��=s-D��_����x{�v����-�H�XZ�")����e� JN?奛�t?�^��5�m��p�(��J_c;���c�γ��ҠG~�{NJD��FN����":C��L�������Bu�AO;Ud��)`Ǥ��\2�T(%��TǠG��tu�W7�����B�pT�,��pB��N*�g���"��a��QY�/Hm�h�{e�C��_W�#��:�9j���h9�PHѕ������\Nox���,�������{�<�����)�2�d� m�"����-��vc>u��J�^�j��^G���^��,�  0n�V�Ce��&sI��飜�C{F�H�3:�U��������v7������F�\�q�:�3�쎅Z��2�u�."�pKFjl.!u�M|�;J�b��W��t��ėI�_ų7\L++��d�CP���>|>�٬�)��$��~e�%���Zq1�n3-7���h�w���_�"�"C^�� ����wn쌠��휸L3��K�`JRل\�L��R,�NV㏋�5>�0m ?�G���1�B~k��OL:!�˨FQu���yf��r^m�R������:j �g<�qV8�����r�:��Z�����g�~�0�k�P����PU�,٨���6};�1�.j�M�r�M��e��'����CDSnaͳ���v�Კ����P;+��tEB�i�@?��(^}q��,m!A��d�X��&j�]�$9�4A�#�i�G���%k��p���`����M����Sb�Dy��ɖ"��.qO�`�lf0�Q���搙����c_�(�¦(�惎�/���s�r
�����v��b��g��P5>[�9+:"[�6�r��)�AHM��Vn{�I�wa����L(ړ��=\��p4��8�u�7�����A��[��'Y/�����s��)l3�>��^�z
;g�RR�׈X@����U���[ w[�~.�zJ`�[#X.=�X&h���Uz����:)B�B<g�_ius�E+�󑔣2%��c�4L�Os$����*d��!8�J��PΕs)�ai�������-s$�U#����FC���7���%�sA�ZEue����󔧣��Z��Yp�E��Ɋw�q�Љ�Э9�y0�=d�h�M��-�V�Yg�V%�v�zGr*U�MiS ��brmw�0.j=�o�@���d��bE���N��o�Ӏ��TY�ǧ	��>����Vd�5}zW��)�y�J���l��RGK��s�_���f�	lew����1�����$	K#���6�'+QW��8�P1L�E�R{V�#����H�"U��c�B����/V*u>,=�؂k�Zu���B�lV��+�8i��)6>F'���%7���|,rB�Ҥ���i�|�;߰�3Ѝ�g�3��4Ғ�����i����۝5-䶒�v׌�����8��d�Y7���:�~f1<8r���u�?�H��)YO�`U.�!,nV�M���e�B$R!M�ۧ��9�A)X��&�	�6���"*�s(GnO+�8b���^� 9���sO�����(:Э���>ɍ.+�@k���J�~��5㒓RZ|�8��X��~�GB�ψz��o���T?�,��k�L���ѣ}b@�6�����5�%�g�^�Z���9�H^p>�\=�W0|�p���b���̫P����)�Dp���by�K@N9|k���"\�\3��H9�^$��
ۋ���!.�t����ε#n~�3<R7����o
u��D�a�uNq������?]��j �6d�I�"x�b���@K�|tk����ޙ����{��51��rf%Sy�ĳ�I��.�T_~ܟ�HA3��{������/�6���)��I��ȉ�'SR��UI��B�m� �#�m����[��AKD!����Kgi-~��,9�qG������=t"}S���W����3�VgCu�(f�Fpפ�Ja��p�1�i�;�.� �>�q�6\?�/�yW�;m�;@s���Zv(�?Q?��j[�0�t"�6W��W/wƂշ/����nz��Ƶ������	gka$�S����s^Ҡ�Y�ʬ��f3Ƌ\EZ��^���3�ܤh?�����|9=���=o��H�Ml9_�_�J�G�Dߥ.�}���[����Uҵ�,�O��t��˟t]�y"W`�}��u��өkJ�d�Ӫ^�H ʅ-����)�wR$�A֭����Q�c��e��β�P@bCU��V�Gx#�C)��G�����9����1{��i�B�9;�m�G��_V���7�z�(�8o�cA�.��~���Ȯ�C-�7H���M����_(�_��ŪF�.p�XN'�2T�b�Q��*���A�o����Z�J�Y׻�1;͗+��l��C��Cq��?y��a)
��O��^�]�+YV;7�q�)��5�?f�t�0	&����@u��LmB����.4���2��3��Qe�Ԗ
a��q�hT����=��t�v�~BP35s�T��S�7�� lSz�we��մ�w�O����k��{�&�b�7���R���dϺh;8m7(2g��:�,[Z��i@c�c#*�X����u&�;�e��F�l&$�K�&�3��r�܍L�OI��32�P�2��K�:8�4Z�U�D���U=���~��A�E�$�,S�h���d��_/���irꪙ��H��N�f�cR�a��P�$��B�,��gh؇�1
�KnInD�B��\����� �mz��� o�9WGg�vҶ�禔���iv� hܡ��#���l^�i�͈�2i��k�R3�##��I�� ��6$�0:��?V'��2Z�(�v�ێ������[,"6T�y����Fd�1A�ʹ�`&�4Nrn���4V.ت2�>�R��y�wT�#���{��ܰS=/<Gf�z�`�����9��K�- ����Q5�����l�����U���>y��Ľ�����__7Y�w[||*ya��(1Y�����}��7s��ɨ�Ф3l{UGPqqA���q� �'�A��r�LN���f��ʠo����W��d7��/+ms�f�0�]ܾ0�n�$�ę�
m�j�mA�=	|E=G<��o���
�v�1r{���ڲ�ӧOg�vk�'��&��1j���e9p��pA�[Xv�N�߷�6�d߁^̐ �zT�Pj9�U�$Ȉ��<k͜WZ�u������Ц��C}�!\vg���4�Τ��>�%XIo�,���?lk�G��ރ �1��M�� �VI�֝��@�Q�SڠE�]���)�3��)S ��u����%s}�<��6�b�Y���,Y�/��b݈!�����ی��%�蓌��pf�	�Dv�u��kw
"1�%�{R}��-㖪�혷�ju�P�*Q���QN�TLZɾHq�� U�6W5G%GXByK�%�e��-�+����${Ǳ,m����Y��)f��u���Fc-!���RjK�s/[���Bpo	^[w�+��&��e��9���C���:��3Hb��5�a��pU;C�%�͌�7���I�n�6Y���z�~k��(�B������t3�RdMP�&��:�W�V-ӌ���s=g�7IzL$Ҟ� R���m�#.3b�ڋ8u(��#M��I��¤�cw[T�;�>w�S1'�_V]`��H���$�Ť�MG����I��=1� 
xBR��U��>p��=�����o�h�����_����D�&/��zY�Ç��0�b��m�S4�m.ɉ"`䶭`O�i�Su�Y�˟!�x��T�p�7k���k�SG�.A�fEk}�W��v!W�; ;z���.q���a���I�����h�ε��n�
��^Ih�u
�&�p�*����ЎޛG�)]��p�ܡ��%�s>�M!׿\u���*f�o�l���Q�`��\``�H7H�b���}�/q��Y��Wٰe�����w��d�ɶ���W�s#h*{�e *QR��o�Ted���P��Z+�:�I��7�T=��X�v$�J5�\̊7��1�Pп��Ү�j.w57�v�~I,l]PB�	R9�
wzW�Y1э�ؙi��Q���r����"@I ��DR�.9����/��V�D�4Q�0b�׋AEh��-�Cr����e��u?�D47��-y���#�F#���MI��Ł,�
>
;k)�d�kuQ���b�9���:3W�����AΟ��j�u���y]6�!?��t�^mRV]��S8ofAK�����n *�GZG׼�yߠ/=�teP~9dZ� aC�p��V�T���#�2ks�a%�-���ڷ�4�=!Xj��U\Bat,~�w�8`��T�A�)'^����;H<i�'����:Uu���
�}4�L��n�6�#~��ٴ�N�E��'�J���7�o�.�ω�q���5*"��-&�'�u�`SuC�������mh?;����޷��#��y������Q�,��ёSX�T���9����� �~���~�5,iB�'��m}6�g|)g�x���$�����7k��'@["��b���W��d~]��U[v��eޚB��Ѵ1�YB�Fw�\>����I�+�z�����]O�����}��!hJIݶ���
�0��bY��$=�'O���=�C�`8b���G�d�6҂�[�:�oJ�n��3��K(Q������E2I�$���6ņ�\�;Y2��yUX�@1_�����?�+�a-3��J�ū?�J���w�m�겁:}g����'�i��kFN*�m���w�����+q�3��W<.$zN@)!� :f��~��/	�:��/6����@yV�A��������$�^��^!�9�w�6qS�dZ���g<�<������7.貰�g�&:�] {:PtP��u[�O~~MG���\��7���,�SGO5���Dƭ��c�����/I��	i���F�J��wJ�����6M^A�\|�Bg�
�kC��\�7�/�o�+���+�-,�XxEH�����L�?[Q ����1z�NZ��6(�ï̗�f������^d��m�b�*��nf��" �)x,ԯ$% N�l̇�_kHB(#U5���F�������Je�{�H��6���z�_`#�G�<!^X�q|�?eDe
ܳ����p��\	ʽk�i�cl���c��!�5��N�j>�_N��5R83jCG�p5Id������z�}�
[kAp��甼e��擃�WF4���2�r���{���Ot�ȥ釠�m�me����ҭ�`� �
^3��F@��9�K����bl�߭�c� �Q�f��[O��ϓ�~l�v�|,. y7�Ȟ�&�*��Ɔ��l��[[=�l�bw�D%��s�2���^��l� Fw-4�.�@�zrʏ��ߒx��7`��kˊ0!�W��k�tˀ ���زv�͹X��w��B9��R5v$����y7夝�j
�F�s��U�vp@F얕Sx�n��;*
���߹��E#�j��V�g�j~��f��V�H�N���T��!H��ė���$=�=7?3�F�zD%�m�J�4�������"�b�К�����С����%f�hD�	p������S95{ח����}��n��\B������i�:\�?�8j8��Y=7Ir��o���7�K�ﬠ�1Q��WP��Ze@����X�[CG��mޤ^�2a,�3M!�0%챳��/�[��	�@�RN�g�q����������K��K��zU��WP�қL������w8/�R�v����^I0����荂���D��Ag*6�ŉa�n�r�.`�qj�������d����A\��`��t���O�#��Zd/v||�P�m�@�޳ʎ�/hz#5���g�.���x��>�'�u�����+5�O�ϫ�a��/T!���D#*b=��?]�V?-�����lE�a}6��[�p<}_�����>&3����5 =3"��h���oLP3�T��{���]�2�;m.rv�z4�Oe�w*�>�#Z�Urb���h�����\ �U�z:�p�����d ��u��P��?��90�^�s�0)��>��ш� ��Hj����x�ft�L�7o�t�����݅t��x�ΩQ�;�V�8#�\�ؒ�D�N^����,�#7���#A��=�o�*���&�˝f
��	�neFs>6�k4e���v�"d�p �S�g1y|��O֯�Z�\I8�-w��	�Xs�3�ڈ��8
�Gp�	�q�,���a�v�"����S�Ld���N�/�X/�D}M�C����I#��r|hz�m����h��G�>?I�(XdO	�����T2�W�ƶ��c�!0�]\(�%��x��_��N5	\t~��>2\�����T!�0�+_�d�`��H2a�4E��ɾ�h �Q&�D/5S��(6K�U�}�D-�W2������޼���yRl���4���a��"sڍ�,�l�����O�J��PR�Z9{�������	Đ`QP���p!�Z���� x�ɹ���`�� H�	���p�Ԟ�^u���ĪO�L��,kh��k="
W�e�$N~��b���F�65�D�cD���qMA����7�D��3����Ӫ h_t(�c+�<>q������vK�" 5F�N@kj"(��K�i	�qrtβ��U�د����{;^���UPM�/-�D"YrF.	�j�����6�j�����{i�*����>IY���)[��iy']�=Cπ�y��
;�����E�y8�����Zt̃x���Ɲ���'Iǚ�׮r��D��Ќ�9y���EY��M*�z�����!W�=:Ŭf����m�q��8�A=�l;���rBr1�]	äP*���7�?���B�lI� w�s�ȹ�7��ʽ����ʡ�փ	�`�ꐅ���J�u�B8��Z���UԹK�%h[},b7��?E�E���tΚ��y���l� ���ky�~d�qK��0�?�%(Y� �N��S��?,v����G��[#��c�ٓ�n"����E?�͗���ڛX����J�uD��C��G�(!�� 2ؼ�+��|8쑭��2�-{�E�j��,�y��m�ǯ�<����w_#�S��筿�/���'��:i���z�D�[RgQ�� �k��~.�ذ?ʽ�w�7ie҄���$�𘧤��b��~a��8������b���֬}��i��kk$�ת)0��l�`%�����ϛ��tټ昣^�}]X7��7aO"�5��~��pV�Z��F�����ZjB��w����T��7��q�+���R&��"�Ep���g�T��\1����6x"���ݤ��E���CZ�B.���cVteF)+m��#lN�~]Zf�e*�� �1D�f���- ��P�������|~����Ad���7��"|�K�ˀO�z����Nh=��jch1�� {��r0dg\c+��|��T!p�=G%��L�{������~�=��J.��r}s~)�ހ�?�C�������c��cv��Y��	�U�n�VF�?&ĜM����tw��>�1Zu���$`�袭?�P<���/��q0�d4 ��ب��|�2܁�X��j�y�ź(/9QM|�v�	+4����Ơ��R��'i@�Hز�8�ǕcYX�=p��ѧ�Ŭ
�$֗��֌7z�/n���G,�#���a��@�Us�g����e�qH�xJ�T���O-�i�!@��4l�/a�&��yI)A���\C��p�B_��R�N�Y�7n���ĈӍ��⒊Mw,�I��B5W�5�n�.������n��u,ҡ�k2\�  �����OL���K��Hfn����e5�iJ�6Of���ٖ�~i]y�k皕��X�e�T�6��j�t�;Pv����L����"��1�xQ*�{w�Ea��\�c���:x�H�ӂ�K~1�\�MpE�CO.E@Ҋf,�M�9�\��po�X}&��Ck�ɥ���� ƕ����b��L�X�Ⱥ̃^�(T/h�뙭51��Kq}}��^8�O�Y6__;?n�΁ju�/m_C�J��l�vo�,T��a  �n)!��f%&�(�<�&4�j0��8�`�w:�7�<�HoOـ�^���Zk�㵫l6�h�0ǎԵb���%ıj�����O�����am]�6����	��������ʿ�tO�_�f�����=b`�b�C��	kTn���h]tX��D	r�Xo.o��� ~�{W�+�W��m��D�f�)"Su�^�>�r����z�_dq���M�i��}��,��u
�f�$�L���;;�����Q'�'M@G����p9m:�P��d<p�8W?:�锶N:Z[�?�*<��&j����"<a۰���(�_\8|ykD�9ʠ�7�W���{��T5��1)�A�w%��@yyOM�$���~w�U�s�(�^���*V�ot2!(�,*��� ���Ϝ%
�Aa��<)�^�J�y�_�OV�V���Z�`L��ԹY�?�jM)c���L��C1`zO(�u3�{�sw�����!fabD�%|[�[��m�L5ּ~��y[���?��M���4m�T`���Ç�_��x+k�y���\:ѯw������7]�v�CS�l��M�S��(��:��D�S���2����D=����PF=�߾|M<��E��s����ӥ��*6M&�Z��mu���U��q߽X���Wi�ή�SX�N��c,��W��^�:�f��ֱ6��G�:dD��|0��b�x��ӯ3�Za�J�<���W5(�<GP�����#�L�K3w;Eߒ)k�0���g�a��gRnlg�L6��k](=��k ks�Ԡ�Jٸ�繴b �D.�CĈMb��X�5�ޏ���<]�Xh�[���p3l�ՕXc[�h�N}�t,F׶TN�D[����"~}Gш9o2���k-<{KŞ��Q�SW���w*��]�NF�=y���~��$�Fs����������xW�l��9�3"]������o�#�D�6�Qy6W��;6U*F٢����6-ť@����)?K�Jcɹ 
� �#1���T�/�'�e�'���E��I��������9ja5v�`C���;R�p�6|��{��fu�|c!�;��rG�����I��8�n޸����P�r���E,ɸ�h�w$���l�;z�Q��i�t�����>����&d���7���K���[���8�5Ia	��_}�`Ӵa�Q�����&�K&�\���SvT���[�
�^XKc�������f4࿩W��}�����0}J��IHH�:��_Y�)�_xz��c&�LIA2�Dz���p-��;<e�%	�D�0�-��yrcS�q����F
 h��=N����67��\�I�u�����6�}6���s�$n�P�������:C
xv�(�S�[�)��@�D��ބQ��R���w�67�Ҋ�@�3'7\f�9�,�J��Rx8�@=�<q�Xa	�東LG��0�м��/�e��Y�3����=��:sG<]@�4=���lkݎ���`-��C	�
�I�g���#���-8D��`Z�"�C�߁�i���p���='�����D47�؃�,U�4��nN��.�:���&2Z>}A�n��+b�nW���P��}=!@nr�n�}����Ez��]J�Jtp9*zթ�
0o��j�����-��j���0�l8ҵ���ǚ&�������;�ڣRU	%��+����ҧ�L��U&M�_	�=G�z��P���6v+@�:e��Ԣ5=����Z«Zcz�0܅�YN��G�	*�@Zi��<$����t���OK��:4��19���A��½� !��Q��-����]�ߔ���cn��X;ɝ���G�m��/�Mbc{��d ��8��h�~��Q��ʸ҆���\���N���bz�)>�ޝ*Y�y�n�H5c��S�&�m���w7*��0�%�k2�l ^��l�`T�сO�Q���)m�@%�4
A��]��d����y{ג)Cd��:��y^����e���U`� %��c��a�y*nO �V#G9����#���e��EJꋙ��"��t�-mW��a%�=*͔��/n�85{�>��/88��*G��ᾅ.0�z7���ݞ����i�b~R50 O�>�R=����e`⯁c�^Jv��54�6��t�I#� 7��rQ��L�Lݗ�:]��nX?d2UȤx�mr�ݜ�y��:q�c�}�a�KSf�����tۂH��a:����5�.���?aש'%P���znq֜�ضgܩjX}g��e�G̠Y��Q\�ve��U}P�h���G#���Z�X9H�h!C��[�:�`F2
�{h"{��<;�hq?4����o�$�I�w��˭�*���`%8N���X��w�s���:����%�
H�-�ɛ
�����l���W�~eUi�L�@�r}dȾ�6�멵|MP`mw�f42�V��8�b{c�Rz�"� R���&(���л#'�s!��|�!�?
~���o	�$���s2����)�}�U,oXV"���,���I�nb��.O�3j�Y+7D5�F�n
�@,�1nm����g��y ���»�Ϲ�8s�t�if;;*��!�B�ʺ�cJ��%	��K�Z[��� 	�M��2s�2�L�i�����M��M0Fz�84�IMWJ���b�(C]�N`����΁j����`S�Bb��[>;�D������Ysl�dW��΍Pӛrt��]��7H�Ń�QL!�Sq/fI�Qg�	2�{':d�T���U;�+s���>���l��R�������\�`2�x3>=��Aq���0�m�0�Ϗ����Q><�1��%�c����E��5Dq��}� �r�kGf�Z��!Jw��<��?�����+�]TJ(��|�!�	���$6yKo1�؉�7~��Ն�M�P+�*]�Π;k7�����!�;��(jV~u�>(ef�:J眫�D�-j�u�#���J��j�*�$NR�F��n��3�n��Ja84#%�����%
}�.�^b�J��`:���X��{,F���
�R����.~a���\M��w�|o���`���=(&�Y&2�jEMŰ=��J��b��m����8]>�Ms�@�;\����6B���@�}\���������|=%�=��*�����(����8�W����]{��ڙV�?�-aGb3i�ۆy��v����ޙ"��3\�u�����Gꪏ�����ΡK�0!_��PL��U}��»�5�M���D�4[���7���>.+�������B	�EJ�}@/h̓f�&7}<A��l��W������ݳ��k��fJ�G���I�^E��x�����c3QX2�t���M
{�޾Ҳ�g��;@A
5C�?��F�M����3�a�Ù�\��c6��+l
����$��B�L�� f���������W1J��~�\N�-��3�qL��v�Ȳr����3�F��uf�4���I��y����% F;@[�L��Y4Un��6*���{d������l��P��Ox���/=IH0�mjq�ң��B�/;�cKC_�o�X��P�X2
�I�K{�ЎA�@�+9.\��4%��� �		G*��>2�*VbA�J�K��?w��qE�B,z��[�3З$��P��uÈ=��fQ�/��w�pܳV��m����.���)%��A��=�U�.���������[Κ������&�s�z]�]���6�OwHs�Hu��dY��:��1)fQ��@
�(��}ߊdH���:�E�?*�$���#"a�ڬ!ۅn���y���d|�l��J^6��G,��B��IYӵ��I�R���0�{�_;�����fib����fnm�v��N�GCh��d1
��>Eg/��$ȝ]���-�FZ;OV����5׻�#�I�Vf�Z̾z�i�i�r��&4�`֡���"�Jz�� �Z����D��,�
��R�e=A�-�@��"�Z�0w`�M�M�f�Ԋ���4�#a���:K��Ю'.��x�� ����9��f���0{�,ʰ����
��F.������g��9�r�W��֏:d!��5�g���T��A�����,y����"T��;�94gHk�L�l�<����Oxg�Y\�C�r8�5�>���z}���+{2n��>,��aҵ�,�h��$�qT���6{�\��@)�|G;Y8t'�� %��i4���O.��5S�;�\�_�^&1�V������=�e���2�3;���{Q��s����1n���c�����Do����{�O�壾,��^S=�s������SH��D��0C�5�TI,����b�aٮ�O3G��s���=�݁���Ṁ��(�#\d�2%$�Vs��-x��j�L��M `&�ݽq��~��}N���S|�R�d� zv�_��E�FZ}��"�]�ƚ@>N���&Q�D���h��.8Y���i���d�-�r&Y	���Ӟ�6��Ad���jG~
�3�]2T�Z�<N��J��=�� �%OIG��(��Z^�f�����D���P��;V���l�y�+���42no�_K�ʼs[�Ff����M�v�GEQ/��j�!��(!��n��,����'��ʏ�]�DP�6��
c+�j܇Zh/���1�O�ƍp]�C��]��_ęm)��Cw��|9$â.������e���[إԖ�{�+�S������A���&�g��f㢏I�H�t��S}�y�9�B�&�;����"�Z�͋>+�X*�Ru�sn@y�*H�9�8+L�'���k�&�^_�s�9t���E#�ϟT|зeo7�m���lM�>�ws|
�>L���01K�dM�1X]9@�:G5%��&f���]�$>p*�E���d!�%��pá7<��d���
Cg�C��m?�������00�[(�#���>�!FĞt+��u �����6�1-���lK��;'"B:u;��z�\����5��{��2��⧺��蠖k�n�^/���_�^��DK��(([ho���+z�~(>q&!�jj�Dȋ�g�<�zbg���!ߔ+n�ܾ1w�"/����'�2���_����i���'����
v"ڈm����l�C�7��ou��MԗZ`��S��I^<��i��q�_ ��k4ͫ��o=��!fN�9���%~�6���1N��ey���$	S$��l��)_�����kD3�Dmt0c���l��\J7���B�=3���,�4%�;c��{YV�+��`1�[5^'��2�e�\A뛡m�����P�x�@���ˉ�w5�tg����g��Y�;0n$�,r}��$��l��[o��sӺ/�-Ɣ<���"�⧵�vΜQ"H���,tk� ����*�w����I��kDRC0��/�1���|��vG+���l�f�9�A�Z��BY7����U��9��/�S�a��<	�[ԣs�/m�/@j�G��6h��u��S5�>K�>?�Z��i�2�`����9^��B�p��M�;:������5���ӹ����F�7���o�!�8zg2$�E���eU�����?��1tH�o}��
�:����W�m򃂋'>@�=�O�z'�'��8��HI�-�ߡN؅@i�_���Bw\Џ�?���Z��Eƽ��?���K��[���
4�� b7����w�hν��\��*�+�=+����H �>s�{�L��/�x� �Y���̊~��aI��a�˙��)��o�[�>��G��]},+I� ���E��QQ�S)�X�"Ct�I2T��{���O�]���޲\�?�/��֏�e ������L�z]��s��xa���S"իl�&@�5(e�k��!��J����s�)U���a�R�"j�`\�T��*GҶ��B��>UՓ4�bCa�I332m�#�^���p�{rW7Q&t�ڈ��V�����QuȉPRnj����g�� OOM�x]Gf�%HIN\`G��FY�_�\ͫ-O7ȥq�2*�8�U�c�!e��������3��L�ؚ�L��2��Ȝ�{*�Nas�ih�	'$�0��ܛ�{���s9đ�a�P<*���f�z{�gf�^N:�٦c,s�}$�1p�­WaB?���)e��0�󡀼���$-V�#`�=��\з�d,mJ>o�N�U�vLc�|G�#*?bԝ#�eӻ���2{��4�(���v�ϴ}���n(e��PF1�MR�>�Y�9]_��t=��bT��q�	p�u�)9J$�~W�Y-(�;��S~�����F���"`�d��'��E�����OQ��V~@�L_	Li�T#�b ���s��L]렏�1�=��n"瑯Bpf��+jW�gځ�6�лhJT����@��G�v��h������E�����I%��	ad�0�t���H��Y�r����:������w7��2juJ��;�Z�.8�̩�ΰa�rR�0��(daq͑h_�~
氒�0Y�W��o˪Ys�e�_8J��'d�h���?��`߈9'�[�̨�3�C���_�n���c�&�TH�R$�>>Q���3�]����c�����F���I[ �B�2�\�r�����rq�]�����1�z�����^6�,c�g���vf�Ǻ��nѺ�j�;����K�=�>V���܀{�D�(�2p�@�g}B��k����tٙ=|Rx�-ܚ�jp�t��	�ŕ:^�_��>�ː<��{Ŝm��5i溳M�c��u�Է`�鷗dbN�u�-���W�e�@��Ҍz�Sw���!-��1���v�<������4�V��r:���D��&�a�V�qt��P��}H4��J�H'f������T55��`IEd�.�!9�=A������=T#OnU*�3�g(�M-QᷝB���.'��7�xo(mD��캑�~��I�2Gd0#lq��&��7���7��Q�	3� ��yL�6��@3�Q~�|�Ia_�dX3P�"e:m����~�#�#[��eu��сW+9�2J�hc�_͖���T.����������d����[�2�˩��Q~�A��}�>5RץI-/R̇&Ԅ�ݲ���ʐ<,�Y\�H�QPۼZ[3g���\�cP|�XG�s݇��^J��?��@�=��]$�(���m[�0_�v	iC�B�|��SF����M�1�M;酕^nž-���}ku�bs�*���M�4�xu��8�!ī��h+�O7�n�ø�S։�*�xo�B��t�c��l��}^&!�@�T��9�%����z���%H�UL׃��΂6Af�6@���n�?� O�Y)I���#X�Ȼ�F0�UR�����P��9�3���3Z�7P{��[�:e�j(K�f
�,m�������:��a�<p<6��. -�`��pz�@�����A+x�̏c,R0n�𢀑�hVz�h~��gs�CV'8�Ly ����%�n��މ�%m�/~@O�6���ޠ�ƞ5��8v�T��p@l�Ka����u������n��4=���R:����kȴ#���o���s�w8ǩ�:���#̯a�I�W�j��z]q����3H�}�r�=�5 ).�:��_��d��Ÿp�B9*	����AO�헸�W��h�R�ʫM�Uo;eycQ�;��q)1ÛB{}��!�MP�u��?��7�Qs�\�Lc����ɭ�r�F$��}�#�_��Ρ�Q޿��_tx���,��4n,ٝ�V��WK2����N2}�$�d��Q�2�4�֨�Z���la�`n���*���h�[R�b�]���c.�x�V�́�J4���f0����%�?'���Ɛ$�����ڞ�)<N����_�w��<�E:�B(�� �᳟�q���%����e4 ܚ���-=�2z7��r��K}ǸZ�9?	�H5x�}�B�%P{����oQ���A>(�0��pL�{���ˍ��5�<z����4��w�m
|&�d' +�3�TЄM	̏��X��X��	^W��0& h@��ݲ^���k���Z[o._V7������v�vц�N<�5�#��S��U}��:��"����,�9vW	��@o�r����=7$��T�/[l64<<�ՊE�����hf�����;��ͷ<p��S�cq�T�!������'FQ�Sm��W�ƶ�rـ����
U�U*�����V/ޥһޓ�&n�l��Ӵ�Vَ{�̉�<��l�9����`:�:�|�̶����l�!��N)Yƿ-����DRo��6�Tz�~0��Ɗ|���{`Ww$���Ǜ�2yW��"�<t�Q��=2�bԎ���^��rr�e���ı�بV���C�-�i���p-k���f��@�T�[� C����AfqW�8�������]v���|�fiG*��O�MK!�<��q؝���&,MO{�p&+;�QcOumYC{g��ђ�t �!��Own׊B�����σ�?��J�V���A���Z�p��X�����Z�%�͵N�{<�!	�2_m_kP*���xpa3�(�����%�����_8
 �C�ԗOe8,�H]���pO	�24��p�+ST��w(�_,��Q���C`j�bc��h��L��F_8/zΓN��wy|���k��f~�wP�����r���Q�,�c0.���f��fT��[ (S�b�=�E��<%�).w��$ �9Sg��P��d2(�����ߢs!?�T���"��ɤ�'؟q��.�9��Gyd��J��}� �C���w�`zy6r�]� �fW�)����l��C�?a�:ĸ��I���`��^!w��Wr��G d{�|�U���p�zH�J�;�"�@v��1��2�B��1���i�7s����$��1��Q��b�/v=x�����oN^��T���Fyvm��n��
�HK%�W���9&T�Ks�rʘ�Iy?�#h��5����n�s��,!�'��}!���7�Z�3d��IK������Aym䅇:upm��f�b����E�c9N&�U����#H/��ٟXr���{W�dr�TԄe�?`�4,��Y��fj��C�4Lv�Ĕ׍�o3=��LgiyGR8I���'�Mu� ��<u��R�|�M]�r����W��I���SjC-rBd)(ɗ�J�E�-��+7`���OH���(�5G� ��n5���(�PW"��Fs�bR,��Wo�"4	���P�.l�oz-��r���SB��ĕH��'ģ^�����G�iӖ�9��)�id��ܚߏ~&ݾ*����"�������$5��?_!=�	�p�����
Fo�|j������>�.�}�8k�T<�t��j��s$��.^
x7��gQ��?F2�F�Y��m��Y��╩C���-���;���1�����>��B(�����ˢ]�L�n�>�3��o#��>8SVa��Qh�m��_1�n �戽�138&^���"�JlV��IC���?eQ��G,�?����"�K��h�P��I|�^�eϫ��|amƺ���Xk@M��g	`k�+��&7o�<���`�X�\�*Tx7�ͩ�����͜�ܙ��>�AW����C_�cw?�p�CǛt�j���:�ƌb���œ]O9U����Zg�߹x/����bd6��FDD,<����_�0ӭ�M-����/�ނ%@��kʹ{��%��J2e�eC}1Lb���wyJ��H��(���N��\+P�سc5^�lD���`����W&��s��o� x��R�
?X���o`�c�!��-<�ff5��7Om�<ܓ��>�� �l�Z@=�N�)�P�t���!)$��C�z���۵�jn��e閇�t��.����G9Ϊ �&j���>k<���2��4U�X�#�>�1�����f���4_})vك}���Df��nU��5_st�e�Ӈ{<�ǥb}e�� (v�Zv�+�ZEm��W3ݪ����F�I���6R[DD��nB���TW����v�=!b��W�̫urm����`m�*cs;mi��2��FAYY�v�R���؝8��`���{d�3���0�e��t%L|2o����j��q��V�E�%��>`�����A^{�Y��Nu�C�!קR%�»�|:�oG�e�� n���͏�@A���h����]�٠�Q$��A�4☟��7gQ����b*��IiBV�=����)[�Dd=y���1�Hf�j�ڟ��Kƺ(�۽�ZP�V l��j^� W?�����N�X�P��T�n{�| ���/���tm���7����f	&�+�m�f��>J�!�}2{�<�إ�'��w�̰�ݖ���W:�q�l����[S�I���A}�YD��pp�{QC������ò�x�V`[&?�Q��T_�;T��Ӧw�CΛjwX=���D-5��G���0���L�RR���X�b��j��H�7��Y�Gc�L��-r�=�͋�|�����4�K��x7΂&��Y�詳$a@Ԡ�%�i��2<�Ʊ���L��@�:л[�옰�.��O�V���DGh�=��5V�P!��D�o@�L���.��*����S�LN�R<�_�
F�8Wz��P����X@K�5��ɧ�s��n��~x��O{�3)��b�M)�UI��m�4�ZZ~W�-��p</ �>�[�	|M9��/e:߻��7��V�����n߲Y&ـ�w�T�3�L��� �M%���� �f�2�n��+���r�Xm���Q9��O��M��� d}�J
�H��S,<*���K4.��:�W����FLָ��֡|��8V^��ab�$Oݯ�<替5ꈥ�4�>'��٪@�ʍO�N6ڦ.���#��jk%���� ����d�(�q�P�3VF��j�f,3�=���!��ɒ��2�~2�=�w�W���ña$��P)u}��Qo/�;�3PŗI���"����;��c�E���jL������l?�5�-`�G�L�aBs��{�+BĦ$�:Ǳ�No;=2��^��AXs�Bs�
����ah�QU!� �S�b��w�2P��h*,K�ߤ��� �ғ^��.�� ���~&����^�H�� �G~��WG����%d����r��Cv�7�}� 7����'�˧�}c�n.��67��F[�F�"���λګ�S�C� }S[:DJ[��X�P<��+u�5�������C���$���0�nl��F��e�8�q�;2+OVB��ݡt����3o"P�Cc�,$�fXs~�gLS�ţ�m)���#�V�ӟo؄ �E�o7�ݭ�Q��4�''Jʱ8���yۧ�,/(�o�J�W��\��'޺O]�ar�k%��^�f������R��]#>_~Q�d�� 3�]��p�dwC`	�d6'Y�(!:X�%hp�B[��8ɣ=�����|�K	��������x�*���m�]���pq.w�Q�u)��6���I���=���2 �c���
�ɓ�Nl ��l��c�{q��!'UV��9$�!BB���EDx�����>��X��\�*�]Wa]Uw�Q8�`</�p�u�L�&�a!�Ch�=愎�j�~*)CE����R]�f��^��m�P�W!Je���?����c�X�'hi���2:���a�"'�S!t�`>N���x�o�LQ�-̺�q E�ʠL�:�a���;N3�U��ɴ��4 gk�:D��W����ܹB��@��&�~ʈ���[���\�8����y>hu�l�~��<.66��B6�ٮ}b��?��k F�0fG|A�� $sJGHvr[Te��6l���w�o��p�T�T[����ہ�5a�����9u�{�G����O�m@J����
(�TZԅ��lb5T4�>���Ex�l�lc�2v�d�wIP��p��쳹O�H_��9��EQC��S�5N'|�[�_���*�޵�HI~R �0�$�n�<uf�pӒ r<��%��#..!�A�[x�����ͧ�ȑ�� ��]|X �W�7G�c��j��Y�V���f%0��+U������)eֻ�~��[�D����d�ޯdV{�m^K�x8:��h���#��0�֧��vD�~ ��Ye&.���i٤|��]vQ�R�0QM����Q��=�Jl Riq��+���v���2 o��=M�|�mMi��
���1!��'1K��I�{�� "Dئ�c�n�⫡ݶ��5<�N���֣vu��N��K���&��©��W�Q-���GQ�Ɲa�TX1_�����H��E�ʵm�1�w�ʰi�J[�������=GM��_�b4��d�>�?"��t��e)���#���2�D'�RV��&̴&��jI��lM8ߔg�������9F1�֞gww~+�t0.M9|�� ݞЧm�z��������J�h[�ј����r~tJ��A@�X�i�V�-һ��HY|������`��:�&�)rcՍ�n�Z��ZJZ��M]yzH���ˈń�ٹ��p���1����ʨ�Z��9�(��8�a���x@���F�#��;�u�W-�.Q��*gŭ���>�"8�䬝�6,�"پa��ذ_��C���#�BZ����iS��a�U#�PğI,s�AK,����6�Ä�X4�>	K�?i�C�Z�!.��x2X��(D �25�\��$>��s����Po^�J��s<���u8b>'���{u�/��/8z^��Jɣ��)�H.걱zҹ����H= �Y�ft!�<𚱤wz]ZJ�ik����7�Q�/�wZӾ$��Qh���	ת��tK}T������XEO��O��k�UCSn�j�b��K����o���f��b:�E���JF���&R�^���O!?�]�#����q��TWIѧ�!����N�g.r�u
�6���	eqDh��LR@;�2��H����C�-S�x���!?g��L��W�9�Uy���'�)�A[Ht�m=#�31�����!Vj���6�_U��ل���$����Y1�5)Rhn"1ߎ�:@��]Y��U{j�u�'�:��
��x^�w�z�v�;������BݎE�pQ�%��v�Z`�=�y�+,�ߖH��	J�䍿�3�?�ȸ��g��+]@hnVD&���j*bd���L��E$�+6�W^8�kr�A����>�k�Z9Ix9�늪�"�
Ӣ��;�S^L���%�Eˎ:Ǻ���ml}����m����>R�r$(߫7�r,hC�_�C�[��v��B�h��V�����;�����t7sT���yoB��I�J���/C֝��*lϔ�_uӐ�g�I�[`�3�9Jد޹ݨ�#�s, s!���c1��W���AZ��3�kc��>i1��`�G��4�1ݘ��S�PΖ~&�<�k��f��Y��̰˖O&j
�?}��Q��cr����*�tq���l�6j�(a�Ư����D�s�A�V�i�Q�9Yl��~��S�fO}t	mfZ���X�FtC48���CC�?�7{O�1h$�+��<2w;��JQ�NA�Z��B�RN����?�$���5���-\�4D�~�I���ɤ����{�(�k��D�-{=9hl2"�-)s:]��K��#="�s�ȑ�'������I�E�q��,���}+"��P���Ӥ��%c A�%�Հ �,��.zfn�~�� ��xt+�S��T�ErxR�:Ց"f����jD�U��`�a���[��ß��e����~	桉�R�E�p���>�߸qפ7�W��
�r�? ��ͳ�c!t=���4ꉹ�*D������8�����㉢e����	,l���&Fr��Y�	�54Y����>����<���h^�e駑0<�0p���A�Zp�`rK��~�Hp� ������@=�i>�̽X3
Joyru�j�D2�ꗎ����B�h�~R���"ͱD�n����brF���&[͓hhA��[,�
�B�|Yۤ?�EuhpL��������ǿ�������؉��t���1ڥ�6���o��b���������+.��S3g�i8d���Uظ�f�5A�2��?�����+ne�#��;���ⅆ�Hh7��L���Lb(� �I$ ��צ*�r��჎|��8J�8�RY�E��w	�Z�P��4L��M-�ж�S�f%�zC�.��@ 
k����Zr��v�S��y1v^}�,�%�[�dY�8�^̤�,�����Kޅ����BN��*H�^�P����S� ����x���4
C��誊��͙7RŃ$er�ge��{ֶsPC\>n@y��P�N��0/*�p�����#�c����(�̷��h$�iM��գ�z���E��������to�����o	����>x�fݱ$�ސ�%G"��W�Ƣ�A�VC}�!��	:���f�צ?��fX���q����ap0u���b⑥n(O���
��e'Hn����.��y�i_�lO����:�uu�� �4�ۘS�C��D_��~���)��TC :۬n.l_�?�l�FTd�=���/]��Y7��ռF���R}]��j�9S�}�n�B�5�lth�}첦�?��@�?��-�o]~v���$qT*�]>��pjG*��S��T��i8���cd�,���4�k�9�����������4�/i	�*���3�a/�d�lE��zJ��?��X�N�8�Bg��^����C�;&L�2Yj�w�o�޻��4HL�$H��X���9�~i=���&�Іd	x��=/��p�b�]��(�u!�.��on�>cyw��g&)�Y2�Q$�����; �#F��5���}{�b̂� ��w���yoej��Yup��ږ<�Q"�$���	��I�,H�R��"�>�V"YO�r�B�ڥ�\���ygVa}��ܔ��;�.�eLZ�)�vh��8Gw4Bmk�� �O�v��	�XV�>�KI�Y��C�'¥����W�[Z,c_[R��"��h?�$��c�qT�����2f�E�;:��tT4Lp�ª�L�cBTT���N�ǽ���_�������V{�!��30���up �����*�����O���r��\�$��\9n��^Y'�_Ta"�8)�ݟ������?�ƃ�-(6��6�� )���\�x��P�
��o��R���n��G�Vxj��]ɤm��%�J����©�e�[�U|���8,E���p������v�[��_3����۸z���g�|���[�����~���#D�;/��syIrS .V"�'�Н�m���� �$�l�� �I����I�rΣM�TX�Y���`���+y��<��o���Ɓfjl��/?/���z)�L���J���x����7�U�������J����b》��֚��J!j&����w��&;�%A�1�܄�#h��\֧��I��5e�^M���d��p��}�EG��`ž��8E�6�@s���7���x��8.x�jjİ?e��|�q�\��0��
����M�?ї_�]1��O�8���z6�E�ǈ���*n51!��`���=("Tv�[;5��82d�*5I���h+
'{{�:�_�����^m�J���)�� �܍�L�!�Y��+ڏ{�3U��Ín�����v����F��Li>���G�i����B������7���)/0���͡���7D*s�on(�M���2w�Kj��-��a gzn$���װ���cH�\ϫ_ZS������Z9�����O<I��O�����z�m3����㲯%~]��VX�WW��5@_3��
���eh.RDO�V1�f����\��%�����#3��"$���ር&�쐇��:ۇ"�N^1��\"a���*~�c\�����~V$S�q��{��7fe]�#*��^�p(I�T�f�
e�q`�)�ձ��-c$03�<
�ٕR���Lp�u7 �]�y2�X�{��<5�U��JǛ^�d~�?F^�{ԴJ�+�J�?���k
���s"_�^�&)9�R3��:4[�	׿��3a;$XY/MI����#�ͬ�&k�o�jsS��O?�T(%�p�����w���"��k���y���e��p)E��� z�:C��S��h9��f;ו(���j`lB웲�'�^Ԫ�=�9��|� ��!�{3��3�Lww%S���N�{����;Ox��7S3M�D@�t�LlP���`�
ԭ�����@��]ÿf]�\F2Ej�ߗ�f��wԺ�}�1��G�,.�<i���a�-�b]dh�K��U��+�;��;�E��v��>����hAz�^,c��SN�/���h+���r2� ����0HqYJC�	|d�cb"�>��5au����s���
��Ƀ�.I��!�.Xr:~X�ܞɥK�nV�0S�=�TXy�FZ��,��btf�ɖb� �V�J��OkMD�
�S�`����ؖ���d�.�c0 �{�
��.*ߍ$�eg���!��9zv�TM�Z@a���* �'q�*����סq/��\������.�&�(1v$N,as���k�X���U}!U�ͱ�R73s]0�?�L������^��U����IA%�����oT�#�A;^�'y
e@�p���s(�	�O�R4��?�5aۚx��Kɰ��q�X6�����/��|�\�����~C=qf��̤�j�����a{ �ɜ�ܫ�o@��R�J���<o5ө�v�@I�_Dz��i�� 5�RUc9�� ���,�'m�0aTg�Oz�^���3ꉜ���_�h�K<RF~R���ӂu�KH�i��)3Eox�XWD�ϟxɔ��t���HJ(�[ȑܗ^;������!O) X9y��.�qv!���{✓9�WI�����d�}a���=�Ġ��s�[1@��rfQ
�k�J� ח�.�.�<n���YL���Ei�^��#I��r@������"�����PtٲyF�`mm��3�8�E�ɂ��H������#��^����\���sP
�����@��T�-�#w����{,�����y���C�{���X�¢EQ(>�r>pf|1[��~���>b��s��p���n]<�1�`�˒;Դ/Q� ���|ё�&a�v:^<�Z�̏�A����|��5n�΀�\W�(�\�$��(�W��쳈�[e������Eo򍖉P�&� ��@�����/La�LN��%������C��b��_'���}����փ�s�����P��Ӓ�Y7qQw�>֢��� ��+����Rh���ϳÿ�;I*D��1.2F�2y
c��+���������;ń��v6+z��B���uP	F`6��](��{mWD_Dl�3��,�sC�w �ily:w3Q0:W�B"e����A:9t����N��E���^HU�lA/�Ȼ����a
(���d��x���w?�k�7�tp�-w���k��֕��\B�>a��tqИ�i�vX�Jy�`d~r����	n^�;MeYc5�O	P�w�����	"�a0C�Ca6jS8C_+m�^����h�/�p�qQd��`q��ڐf�1^��½�E��3��*i��D�x��ĭ� џ�9���qڸ����o /~��w}c�S�Q	�k�ؐ=�*�d�E��y*�TB��F�.Z�������V��H�2�,�ovP�1�C�I��Egժb���y�덞���K{�������Ø�)ް�H��\�ю$�� +�M�g��wnZ9T�Lfq�#H5����Q���\�Y|�NҼE^������v~�z����M������S���/'7F��b̨��lJ�DrZ�D齜��8�$�}�y���+X)�5�vC?�S�!��I�`����a7�^ �h����ƚ���� 2-}�xK�d����5r3���j��D �ڀ���ڲk�*��]D��^
y~{��/<�1`cVC�Q�OJ�r��>� �3R�A�U�9����UWj�D<��۸P%|l��(5xe&��\�UU5D16���	_�BuHH�B�S��#����f&��8ZR���XYu�}m'q ��*_g��L�W��QW�CL��.�B-�e,�jM��.�m;��W4�©@J���b�4"{���*5oa�2���̎II���7_��\;�)(�j"�_�W[� �7A�Ď�֏�;׭��b,�7�0�̱@md`�\jJ���@'�ʀR���0��WC�N NY���x��2j(U�2�m؞��]��3aY[��f{�����K	PP�R�h�d��~_4��2i��K��7xxVk/�.xؐ�zy�o���Qߧ-ψ��>��g68�.��d����K"4Li��8�\l����)c��?�c{y!y��c&*_�Q��j�-��_��7Rd�~<۞f�L��`��}��gz��f��Y�G� U���h�>h6"�(�a}p����Խ1'�S4t����2����5hV��#L[�3����X��հ)�x�����;���|��q�r���4$*���m��@�|(4�]�lֹAk9�GqF��3�jUL����q��h�ϖa6?u]u&@K�����q��s����:�H�?��sYT���[�?}j�̶�Mᒕ��I�B�K=�7�s���f�Oݮ���
�cH/��roQ1(�ҹG�I�%��l�"��ҷא��P�SZ*�졣�-#L��W��%���)đ\�%���>���5Nьx�;Ui�m��f�I��3'ݙ�ݣ1�z�ޟ0*%r�*�<Q�35f�H��"X"ŘW�pk�5�DvQgֳ�2���IV5>�k׵B��v��'�9��ԅ��+_�Y��x��T&��se?�8ʥX~�-��[�e8�2!���e\����TA����q�ڕmz�tG?@<>�Ҧ&L��,�������e�K�R����\:�b�qJ��5�qf%ĩ�<�s�ӥY�IKB���=��M(�}���ɍ��OUz��?W��s��2���-VӼ�;�!H !�R�x?&�g�)����=��g����U_�C�Kk���U���GL�d�2�7�6ɪ�������M�K�����b3o�Wf��J�͏��,�<�����Y_��r��Ϋ��>U�+�l�줤9�DP]�~��{E7s�/-y>�����w��@�d�f�AU��w#�@�g.�N������f�������Od�p��?~��s�'{�
�Wڛ�F��r2��c������GI�ߨ�2���7`��	�{���tZ���j��U|�׆��6�����l�.�6�� �F�o�Cv�w �3?A��� 	�����4)1"c��H��>R�̑`�M�v�9f���;�*��P��LG����x��Wg*v��
ǭs�Cl�.��>B#�i�]�/����0?_����]�\���P�B�I`Ag�57��h�7��u[����)��j��d5��P�I�5XKp�;eKl��'sE��dQ�x^�?�n���M��ql�5'p�pݫ�v���^�0dX�O�&��;�o�G�\#լ��:4-���S�i�b6ɻ�Бa&܂��q�4�ī,bu�\�+���g�}D]�n���7���ս�
�E��x��k���{��/�����u�Sc�h5H�i���?�pe�����Ԏ�e���5�ci�W�3'�u�!T�Ku�"���Z�@�@~�D��Nh�N)�)lL�$S�!>�<A�6h�x��psި��`��2��QW�����������q��|;��IN;g���:7u�R�'3�������(됏�"�
�rf �Q8e�ISFCuj�}	I�g�0�����I�;)�\��[0�6 ����w��=̹���IL�4(�oS�p�?.����K�w4y`��]7��B��8�Z��+r[IGi1�=9�*g^t|��Aj�H�i�ʻ��?�S*��5�a��r�kn��Fwm
dDˑ'_u%,�bz|"�h�����&vʢH�j�RK���L������o�T՛'��ꛩ����,�ߎ�4_�Iz1�L���w+a�F�AQ@���R���_Zt�l�~UX����O�c09 �@ɴ[�=<*��2W}=�PĮ/(�C.�sJ@pS=}$��u���]q�g���+��QÌG�\��5�P���;D����9��+Őm.�A6��J��R�ivf��UuJ��z�����ө�B�1o�6Ϡ[��W�8/8����U��#������:�~c�?U5������ű�?�4|�Qgevxݖ�*��EæM�=��\���(��jp�왝�QOø
Bq�Z=Ar"�om�T7BKt�$��L�.�§^�#ӛ�+K�;Pƍo�X�3�������_�ܛF'߁:-6_�$���\dG'��mh��pxJ%坖���ә�����,�����d3����#4���J�.A�a݃�m��8?�7��m�1}�k��\��^QV�~e�a3pX�}��˘��}�ʕ�o!�<��9�0N��b;8?���ǶqG������;�����٪�n��[��8�Rb�1�I�'���D 7�����~���S�L���oS���iI�=�U�򊟼�e!�1_�3^��+r��R;��|���% R�*A1('��Q�O �3�J`�q�46A1pj��@��gw�Bo���X����>�*D�ZP�9-�Ҡ-ܱ�e�y�Yp���&.s4_�(�U���>�p��`�;sjՊvr�sK�'!<o��S՘)�,��E$E��EH�$6D.I��}q]ބ���F�9�7|Lč�@�ܥs�0����>}@I���_�m��q�<�G8�Vdޗ=Q0	z�^�MF��0���i�L�E��A	q�x�ۭ6$��g��dʻ;�u�A�͜۲�&D?&�)A��y^���I�С����b��D�k��˯��=t�����:r����@���'���}� ���ƛ��T�X��w]�o�F��/7o��yKݳ^�h0�jvau٦����r�c/�!Ul��K���ֶ4z.JW0��
~�!o�eQ��A�#ᩒ�x�������Lr� ��B����>��cq�K�kޝ��d���m��O{W�\��!:a���"�Ax�"'��.���G�+�ء���`,|كҺ��4����?6L�\c�����5l=�ţ7��$km��-bM���x�@�̊��F�v��P��5}�=�Ĕ�-ţ��.5�����M_�nO�ތ'�S4��$���%�7�����p.IB7:o7��h�a4�i��*�ӏӨ��4P�"��1+�e��ι���X/�K/�>xC��Wx�����C�����a"UTo�\}���x��|���Kp	t��Ǿ�"up歡���$��n�ԣ��O�ٞ��Y�7�!v�����_�>4��-�M��]w�D�?�_&B� ���h����R�XH�3%7�ce�wE��P���w�Ff���M۪k
�3�����Ae������v���y8?<S�s)JR9����j4;��s�PJ�*���F��/c�9��E]�!$��2�(�9ʲ��n�"h�X;�h����|�؁e����G����\Zh��Z��|�S�+��h	�@eŽL��,-��Nק��h��g��'u�^�,x#^Ӎ���&�8q��U}̔�"��c)�=�X�Ӯ���_5y��@M>0��ۨ����I�;��Z�o��rS�m�S]tY'O�{�EN6*`�+�L��2X���v�h�Q���`K�	�������/� �ٛ�%�ڡ�g��B�n��$�yς��`��#��i��K�P�F(���89y<`���<��2�B�-���P�����<�4�����|��ݫ�t�6�v�`����ƫ���L��d陽�� �`�T.�u���4�7��)�Qg�6��~h5wwW�#!�눝u�H� k)zO̩h�?����_�N	jQ�ͅq�C����W�*Q��t]�B�#}̈�}�¥L2&aKGȡ�����������-���z���W�X;��f�iO���R��/c5���Hq�G�}�RL3�m0���e(�} z���A��Sr��c^$I򔿧�3�E��[P��̯)�:��r$`�I�*��Fs�W�g9;���~�a���\��W�$.�Ǜ�2P�$O�.��|�[��6ׂ�5 M�2�?��1������)�7H-����u+�3��sV@ś܂�#~��`:��)�M�(�D�ߟZ�{Q3y}R�s����HI��߹�S�t�Q��2V����<}��=n;6����m�`%���~'Cina�\��M�h�dY� ��^<���R*�9�������׾^`t�)s��y�_ԨV 7U�U���bPT�5$��
�%���*�~s��W	{V{���3~��� ��d&�x�p���ܕ���y���bB�#�2�w�w��j j��[u������f�B����g�@���]���*����Ci\�>��,�f$w�0s��	I�oL��J���s�� �7�$���������q�g��a!������%\2��N�Za�s]� ���;���;I�[B��u�=��ln�+�f�B�'��o�"����M9S�2�Jn���e�g��oi�N;dI��{�؏7���l2�N��lZIO�IE��	f���#���F+�{���y�}�"+��4�I�N\1i
�'h�����"0�3�	Z|�t�=C$�b� �Kʂ��@ʅ���sczwy���։����TD�#>�s�+��/���9��г+��ڴ�]}�����ul�4��Oх�aSx���hk��=�+T��jO���y�	f'��s�T��Gm�8��|غ�v��;�"���ů	��8���ڟ�)f'�w��R�r��?y19ݥ�f��V���^�/�н�}�^��Z�����d=���fe�t�W2`�7bt�i�d�WU��$��o�.(}�]���j]�������||2�R��G���,^�6p�a�\|`�o�ƌ.f��.�PԁXb[Li���O�#����9_Wp�m�\�B��O����b���h��;��|�M��S�O�B�����#��˒ ����7ɩ�௿m hKxq��)1茟�}b�O1�:7wA���eD����><_R/70ٔ6���q��%�"-�#ԶMI	�*����ɖf��z�'�+��W>ZG�+�I~G�����|�c!T{�
t�w2�:rFmR�Bb)��W�Ŋ�A�$���16�l��]�
�����۳8{	�Sю�m}������pCpW�e�ai�Y�75�����5�-"�w��At����J��HQ����vm�߬�,6ׁ�o8��B�t�g� 5�t\�Z����mۋN%�Z\��H��l�}M��؆�f�ouq1����,�;g�I���;aSsx��LR�K���K�65o����j�W��'���*zI�jJ� W�rY�{x��F� �8�Kz������Z �bw��H# vfr��,�s��>��L�@ٿeB�]��'��k���7C{�
>k����Cm
xG�����Ms��eEa#��*��в�z��L����~�������$�%�?�\���-q�@JO��Sl�e��me?�	���y騐_-A�u�,�N�K+=�����j�f�WU�v�P5�ca�K�����ha �D�j*k��t�$E_����n���uK��>|Ǟ�1q��;0䙹H�#כ{w��]�G��κd�[��O��h���@`�ᎉ�%�7m�dnO�+1�����^�8e�ݙ��d5c�V���C7��`7x�fǅ����k�L�F�d������k���B!.�0�X_�uW�':��s�VATr�v�,yA�h�Z}׏�$��g�K*;q�B7N·�$��s�׽�m)�O��d�m��xƝ6��eqt"H!oLhU�$����\�8�Mc�ϙ��{w_/K��)��r��
��#B����'(_��B�|��ahQ*F���6Ϭ�����h)v`u�~�.׍ie��:C���XaK�=�*`/d��(8�T������g���Ff��"�D�|�=(e��	�-�:0�X���1IW��ܽ�^�^�V���X���gX��$(�����R�d{�k�6h/�8�����h��Vo[|�}�5}�P����V�A0��a���o��q�B�Ѹ:�i��O?͘�* �h���ʙ|���I�������u�5�(����W��"�� �	�u����j�77��[��x\���K҇��##�$�*.���eϳ-�n�gl`&��eGv�jD��������#�MR�NA�)R(���,��:�<�QS�2Hg0oՍ���Wws]E�y�(f̵���`���o6���5�(��#���������E�4M��2I��[ r&�ɥ�:�0}�q��ì�-���`�Z.?�}��d��M%����h*ms�i7_�a��d�6�LTڭ�ć'W��p��:!%k����MF����"�����X�}gL��?��=���ME>G��0���+�e�/�K0�	�� � ���3��=>-0j!�=�uOi$Ĵ�=��jx���6>�	�/M�S��l��[f�]V.���@�c��q1�o����]��?���m�ċ���ћ���0U�n|����ģ�6FsN��j�\܃wEI��v��D��R��� ��̛7�G��R��3r������w"J�v�����=l�J�����#�Y:�TD�������bbb�Q>EJtL6L���(I�zq'g>_����(���P�'23��ՂX��u>_tp�'�)_�E}�r�7��0��udZ���6�� ��7�����\?��,��I����/6p�A��Ӷp�~B�)�ӿ�+�0Ar������B��4
��,����_�����x��6hؖ�FD���j����O�.���D11�{n�oWK�!�|^V��J�&��Q\�'�Z�N�L����)�:��k�1F��Y�I�����,Q������b���O d7�����f����x�mZ;��GX=���3t����U���t�ۋb���ڇ�Ԣ�;��gx�:�8	`�D��2�)��Q�m�W �|:�������٪�{z��KQq��ĩ�����ވ�s����Tb1�{=TV�g�g�H5�]c@*����yY���� �)׮����!�q;r�,w��?'�X�u��#�|��N�ߪ<E��ǿ��	��f����8���?|����W�]�"3�r�%���7\�uE�iةۛ�}�i�u]UC?�K�Ͳ�� /HL�
^}��2x2���BxE��b�ϟ/z��+r\��O2Ux@ab�e�W�!�-j\��T<"�D�K�-AV����tqF2����QP. �X��.����ʫE�ݒ�
�Ԕ�{q���*�!fs�Qۻ
#�X��g��Ň����E_�.1��f� s(������y\�=\��b4]bY'Sx�����M�9~��4Op�>�{�� �]�P'Hĥ���%aM3i�o}�G_��]iE��[�~�G��d2�"��6�sJ���=�PizS�I���ZPLPb}{�3���d�mx���+��}AmJ���#.�fM��sʮ�~ |2�2�����vf���Ѿ��~��nt/��L�Ϧi���t��T�g��F�����賮sa=����kH�{>��`��#Y�$�<������&y����Ex3��#�>�Ni���������n�H",��`�7�}(����/;���g��7�������'�#�b�]��E�Ƶ�4/yK.����+apGSҐ6���,���dwa2�p�1���(V����mC}�.0��1K�F��U&��r���u��s�)N4�!��M�Ҩz��5'ľ��ҹ��h_����"n�i�3R��Dz��8*d�)�.7Z��,�X���2Ѹ�Wl��SHTV�� ���0GU@#������a&D�(�C~��Cv�9�s��%�T��a:zw@�<���T�)YFK�f�O�#��q�]��3�b������C�#-c����J:Nn`��л<]y�7�ʚkBJe}�>���PzX��(��b����q�=&R��Ӹ$cۛnK�K�كa�
%^�X?�pO<�]��0��R��bP��B�I�FAM��C+PS��|�S JWL��Di�n�N�w�j=�`���.G#s,rW�GM�\CB>��N��z6K����aT�O�n����jc|�#���f���b�.6�챵/>�1�'ܬnu2ɕ|H��,�����ɛαxu�}X�t�_�X;��,{��,���L����V��d�n!i��k� �h�m�kŃ�+X�:�F�F��~��~�5��F��eEz��l�@�r�QAJ��Z�mH&�Ӟ�^0��w"�s�Xpq85�zՌ�e�(,�z�	��p\��|Mf3L٤�t�J�mO��9�YAPR,��[�ù"9�j��!r$|_Vp�vH����\�f��$@�c� �Ys_�-f-����qS���yP!�{@�_�ւ:\%�8���Y�bRJ}�F9/����<D)�eS��!�o;��������41TH��_�e�����//�v�A�u�'��h��.�A��� p�l�p}�7�Q�{<~C����#�F������7�Y�*�*C�p���L�>{~�W-���.�F��3��ɥ�}��q�=D�C:���+7Y`��
g���X_��<�(zSH�8|�G"�\�SS����_����Vu�+ʒk{�a�u<γ�9�����f<��G'!�1{2�|)�|���ȑo�
�����Yl:G
��6��T˨��bN���xf��m���]~������O�!���-���/xk44�o�T�տ&xI�mg���%>u`txy_��j�����3ڣ4�\�x�!X�f-���8�FQ.�'�Ee��~��sF�UH,�j���4���D�v�������%|�B=�\��K�uҵx�	T���jgk�u�F��_���?h��q�а6�~Q��V
�@�X����ZFu�
�/2ӥ�W�R��+yղE�"�,E�b�ۜ!k2��zD_��[)�ƒ����,	�Zf�;�0�?�)[�a�P��>��R�
���p����C�m��q�6 �EŴ9��u�B�D4��3B=���<�aJ�m3�q���nr(p@*�0�V�(k�bMKQ�K�����Gz5����e��̲ZV��������D�1�9�b��x\���S�Vp�'yK���<�+7��r~�PQ�5�
�{�	�}�mo����z/��0])׍�q*T�����?�M�xڳ�7B�k_�z^W�Wag�ѕ㫁����zU֝3Bee���7f'Z��x_�_=<A`Z�M>sjaXL���D2p <���vk
*��A74��q�b�[�5sL����U˟�R�U/������E���XH��݆~jMIID�}��-i�g��m����J�6e��"�ݯ@��������	_�I������!˂��F�Bx�P7H�
)Y�Vx���3ڒ����h�M<5�����M���.�X{ٸ�ߚ&��٤�Ͱ�����.��]�T����X��[��Q()������]v�p�'1�1���!MQ�p��	xw�c�h�F�h�����Z���izsZ�t�C��9�)�'��]A�K��w���j!\�)�C��Bd�X1��Ҩ�e+��?����ʲ[��?)2x���������b8W�������n���7�8U���ۉ��s$,�k{ߥ|��H8��?�h#��?֚~�\�%Q|,lVxhH����Fd���cw�/�k*�sBTTr]$�����D�A�2ϕ��2�p��M����1h?�����|"G�2)7A�K°������Ft��pe�@[�DD&��sοE$V���E�>#��K(fL"Vo  b�ȩN��@����j�h�;':����vC� �#�'\�~f̱��i@�1m�m������飛�So8��q�C-zx:o�>{k������é��k�	fIJ~��&�	ĩV��>YBa#�fř!Iu�����B�߿\�~yx�+g�l(q<�8�`��=�[X���.���O]B�:m�dy$r*�Y��
�'E��J�1Q�	Z��x�M��� }�
��v��[��;�i����.��;�0�Q�N��]��_Z����NĕK#��
��F����߆�ǣ����ݑ(�/�'(��E,������/n� �Ix�^K�&dp�~~�j�ͤ���{�W��ƌ΄rP��оL��u�.L)vq�߃���D�i��׿���(���u��N;'"";9C![7��N)}�Z-a��m�hv��,�D'������|2߃�Z�c�7C�(S;M���z���I�v�q(�"���`&�Q�}�GQ�|�7�"�F�=]��[�ގ���슛;Gx�����W�饫э��[.	e���FAߪ�M��&{r��=�r�yT�t�HH��ۭ�Z��{}_d�VH_M����|_��NdP;�F�& :g7+��hK�kF�������8`��Q��IB�,d���e�����[��Κ��1������ ��TV4f9ߢ��������g����2�H�q�K������T+�|T��Z��@�ti�N���B���7��(P�`W�\�fy!��fj>:L�g�7�}�2׋1V�����fZ����˅�G�{Uvi����������?@��d�M�c|?��y0�����,�H`�r}��F����L�r���~�&D�E�:�ه+��� ���/B���Z����̸�f�@�cSĩ��	g����ﳑ�z�	.ե$�Z�/�g�<�)�=;,������B��NY�W�%�5'��T��@���L>���1��a����t��n��Er�{�3�#*[B�@>��e3A���1F~�)�@�"�[���EҾ���B�/��� ��~�/Ҍ�A7*R郁.����oG�cL~,Fa�X<�����eY�,���'n�||0�!�c��^v�w�>��W��u����o���AШ�"�f4���he� o�mn�[�p`������h��w�U�e�f{8L�[&I}�k`n�7�$#�J�Zg6�����^b���c�k\�%쾨-6H�aC�<�t��7��q �va)P��"Q�y�MM���(����j��WI���}��ۣ���-K+�eg1���_#�Q7��`��5{);���=�R�K�d� ��i���S�t�� ��4>��'@��~�E!!��ĸ�I\�7�9��hJ�l���$Se���Kt�GM?����R ə�wo�X�~�.�P�ʖI����}\_�7�b��9�oؾ�F�Uf�ے�tCf+�xҌ<�v���B�ea�S�9���Q؃���(N�-�����=[����M�Mn'y�y��;�@ ��%��!>�[��P"��p�xn$ ��V����|���D��b�ʯR�kZ��q�`k��^��1P9H ��$�����q�cE��#Q.��c�$t>��W��F�OeVL5}ﴦ'�AЩN"��(�Y��_)�:'��f�~T��Nr��Ff�yd���c�(֋y>�I`��8�	R˞IoO�E��*R�z�`��@j��>/���2Ο-7��2u�i@�]���O^��|�;�����(lŸY��pҡJ0��#y5�����^]/ەzhh'ޥ���{�Ϗ��4��A{[��pI9���b����N��,����
?4�z���L���`�xV����и�$�뇐���8��X��ϊa{mFſ�� D3�f?b,�&�J"��J�>pl��#�&���!c0�x�	��H��I腐��/f�����i�2+X �6�R�V���*!�_��\6��_���
�	�9?���K;�Ⱦ��w�F�Q�1B}��:��T�����}�����ղGц����rcQ�r��ĺ�p����E���-�(l���}=�FG\�\a�|�qf� d5u�_z���GxƘC�}PU&��K���U'� �?�3@��,��{{Bߨs�-C��xJ'r������	S�es��@�3Q[��ĖMd:��v-.O�Kq���w_XO�i/�����a�n�)E�u�4�W�P������g�h=�/��@Y�������^TvEp{����)]}��6�T����@�V5˄��f}	H�a���qۺ�e�FerV�OD�7x��EXXn��'7O��M�S��R��8�����{�և�9$��Jr�>�px�iE?�Y!�_W�l�[{���r]V!�T�3F��������`H�&�$�W���Z��D	=�Z	{��}@e� �V���tVr���F8�'i��N�k��XY!���Fɇ����`�L�w'���[m-J��g���a��.I�Y�o�r0Xq��èz�?M�W���'���s���Y�Y����B��te�%��hF�����՛�#���8����F�����o`T៦�LC�=II/���\+s,�8����#ͫ C0�fl?u�kz�&�~%ep�bPP��>6���"xb����V�O�j�fU�Q�^Z�r9q\O���U�+q1f���p�K,���R�yY+��p���?���?�Q�GN�,������.^�0��E���`i�d�p���ȁVq���$G[�ĸd���J?Զ=�7R� /�y�c�T����Kݹ`�v�-p?m��S>��9ԫ/��==��2�~@�J�7ۖ8��X��dZ�as�̰ΒGv6�C��"�;$�|���r��p��<ժӆ
!�t��5�[ܞesr�ڎ_I_���3m��r��M�R�A7yDS_�ۤM����R�1*��PG&l��g�Al�GO�9i��ܙގZK`��˵6�M� �7 Ǜ�T��g�y�nv�� U�:0���>��0�hL�h�����gq��Z+#����� O�n�'~�:x�����+Hg����L
��a�qGv��I&pp�\�Z'm,���t��̡���ByͧG~��181�49Lh�DGPoi*�^�����Z	���넭�_$�JB����L©���S�R�%�����נ{%z:#�r	p�����^���@�CD(���u�ǥ�YD��c�\dݥ��v�<��x1l�i�.����ϡ�"�~��+����X�k4g+�=o���=�x���}���?�}_�V;Ā��w��Z�Q�yn�j���τ�	D�A��Z`�j>2TP�yZ=�5�vLp�`�<�a�Z���Y�V,*��n1��ȍg �����~W����t����6Ȥ�;'S��o勊c�7@p�Ѷ��t�H�M��V�����+�}v_�F�	ea�y�`�<���jF��v�Z�.�L���b
ǿ�*���4D�^��!�$	��Շ�g�Y���7	T���W��%Ȫ#D^��C��v9x��$a$���l�n*��8�\<���r�.���W8���{��VHގ\���3�p:�<"O�1�g����:��la����n];
+H�킹0��F��ˮ�=�.ģ��HjDM�4�|�"��#��Y�Rĭ;�/BJ������+s�+E]��i��!:��W��i�C��A��&**:m�~��%�J�R��@���`��f����v/�hj��4���c<�������&�^��$��7�Lo�k>��Kb�و���i��il�SeҴ-s��]��!�?lR�u��@����#��}\��n5�T��j�\0^4��.�k�K3F%�0�Mf+aN�����NzB�P�v{��E�>#��[��]��fB���rt��w��z�$K�b��^�._��Y�=�3�*n���w��@T�ȑ	�	����*3U��E�9F��B5iZևX��y�@��`���*A��S��K�n�Qq��`��E��IE��3,�(� =�7?̶J�=��4$s������><N�����'��b(J<4��@�sF|�-����x;+Sn�D���d�\���ݿ�^�u�3�Q� �����j��B�#�r@��4ܸywRˋ:<T�8c���U	���ꅖ_K�f�V[��{c�&���G�֙ԛ^5�f tV���2j%ֶĐ{��HZ:��=gwe}�є_nC��$�>�%s�A��k��Vd 6 Dj0.N�HW�p�%�!�� �$�s�(O��X��PLrY�*���.o�<i�s�����;Q2� \��kN�N]m��˂x�,��t����uȁx��-�I<S�%��V�h��u~ZPv�g�bb�5˒>�R���ġ�|�o�/�<rg�l�V7�r$��<��S�jr�7����z�6�J�/]�{č,�.��7�-���=�@k�c�3������z/n�G�+�WM)��kmI�b��7���c��c;�Ͻ�����خ��*W�-�@ 0Ч�������4���co�e�n�� ע3[=p�UC��6�@�Ϟ,��(��am0�1N�t���X���˻a���O�J����/z�ңS"�X��ߢ%�ҥ���Ȍ�8��M�J�QL��HS�G����{>N�0#AY��9�p#=JU.�ߋ9��m��l�(+�M �g��l�~��u$�&I|��'���vC�L4w��?��Z@�܎�{r�I���Qԁ����`m=����@��^U��Po���i��~a>P���mD�4�ׂu�C��	i�X�k]%kΫ����C�F��Zu�b��;��U%�e�$�T���4�ub�B�q�xJ�ؖ�~1��"����:�c�E�Bsr���@�F�z�E����#*�+(�mh�k�����cR ë&�*�H�ll�ء�����W�@���yn�������`u�z���`�`;�`��=((�atv	شf�Xz�H��C2ْ��|���\ƆO��G�6)��\�Zv�(��ѪY瀶mX5����
��߹X���UQBD�d�Gz�}�fjH�B����I�DSI�7h6�J;�<c��=h����QO/vzz}%���A9s"{ g��Ɂ%U�����W�?�{���]*0,�4�kh�y�����^v7M���[C)��<�7o.$,éG>��z�!)$��9�L��
S�D��EaL=�A�j͘�/��d���5jTu��lOT쨯�D_`
�4כ��El=�
��c{��ܣFPM��Z��;+��hi� �)����.�Do�;�ڎX�����V�C	����$������v�i:-*�������ɥ�_y;�4�µ���&��s�n�^�]��gd,��1��PN��.�!d\��Ct��қ�B�D�P���?0������i��A��n�U�o<V�{���H�SN�y5E�V��[I6����#��e�ÿ�/����A,^��w��i'�'�_��W�0�֗A�@;��մ��W�uj���+��T�Dr���d��H�������ul�播��=��1-�U�Ȇ �s֡��<W�/���
��J�>~ҶV�����f�!j��:(�|v��y1?%P���F�T� �u#��A��0\��B&�I��7�,����>�*N�U-"	G�&�Bor��U�>�rE����[�������0vN O�Y\��>?�g|�m�]F��WҔM0��(�})�>�T"Z	xs 9$�r�E�����~�\7����<�l�M���⾿j�sx� �DD�aV~�tH��@�S^��7�R�6�Gk�8��p/D໮ʪ�Y�p@0�@�&*�y`Fh)���E!�8�>�l0"0A��G�MP���
?�Bok�֢	���m�Ƙ��Rz��!]��U|S-��bg�=�9n>*��X)@s�w&�:��m7rt��=<�:�z$8�AA��g�s�oȸ�hJ��+��?s��@|ɷ�ߵ��B�����׾)����n�X"{T��S�Pz��E�e��xu�9�)�0�Vܙ_k���$}��?��~.�E���.��mi����UF��A��T�{;azALܱ�nCo/�/L�N�J�I ������������*�w�24���L��2�����89�f#������l��t=���gƶ�O��f �l��V��c�&�M|�1H�\�&����;�hB�� �a��a��f4�|7����d���a��:~X�����iM����)������'۱���H뼙�V���|��c[�(`�m��fӱ�YcvJ��Bя�Bg�(
�X#�[�K[��O�peչMA޴q*�k`=��8F�Y2B�a���=0����=��G:a�a�� )H靤�Q@����̓_o�,�GF��<��#��*q���7�P��K�����!ն:�+��ZZ���#D��ZLъ�C�Z��b*��<	���l�C� nA\6$�_�C�t=�������t�t�3� @�G�^�-���J~R�)�G�~F�{���1�e�3G�4ABy��h�Gbg+�䊕��#�5��D������&�Z���Md�����p�A��^�w^w��N8��D���ˉ��Q1A+�ǝ��!��@&@��`y��n��Ȭ̳�7r׷�����c_����γ��J�R�����a�7��n�����4�l��(LY�~-�<�co0�< ��q��^d:�61���~c�!�)@��L��N�����S���w?G��ilh������`0h�*ܢH�e���ΰ\�QH��]��4��L:e>�|[>���_fH�慌�l����  Ȉ�?V�	t��y>h=NvB�ŭ͆7��L���ӗ�p�[�r�ĺ�jb�!�lN�&�c�:hk�.ez������Se����D��] �꺗���ܜ�m#��`��]R�a?$��b:��n�2��-%i��ai���s���Mه#S2;��ٵ�^GS����3�7;7�D`o!b�xz������y����W9 lX�A�.AJ������{7�z�M�߹��oc޵��Ga ����V�$ȇ�/Z{�v���4_����.D��,�2�OJ�����l���P�P��((i�v����+�v�S?���V�%°U��V����k�o �(�G���;x<���Ѐ
���8�:fL�,5��~�:^�S6��s�Ng{�T�`�{�d�5�C��1�PkՒ�X��&�!�}���҆Fh�9�Q�Nm�_�J ݱ��$�hu�GC���-�-��B�r�=/�|�����G��a����;��!�@�U����M��#��z=O�[t\6{��,ש�
'�!t-`H��ם��U��Y� ��#���e����ʪH�Ӆ4$�tmU�	VV��%�걤�םE��M�S
��H����b�襶�l�2��.�.�fc,�np����,]�2�+�Ĝ����.W��`��v�<R�Kl��g��w<.�4|���k���άP7*��;Z;��]�T�p�q��!�󔷈�6�-��� �7 B"ƕA!��q�ŵ�<��+��ê}�?pbY�YJ]�������%{�2��j�*U�"����h�M�3�τ
eC���ۚ�DQŶ���:4$���J=K��vY�̊WŲ`r���/6�w�y��t	l�,ɱ���zL�������q�4*���؛���,��
W5��xtPN6���6����؊���Q�Wi��ڞl�Je��n��T���d��~�,hvxy�{���o��dGb�}PO�F O�-Wל�s�0n�'~u	G�]�
��4���-T5��:)0�!T�[V�ė����ܑ1+�
�r(,mi9�Y�T1^	�b�]��8L:��[8���(�vd+y>��ҟrve_,Sc�3��#^���wt�TpA:%Zi�A,�����	�l����m\#+�@_��6ɖ��PT�%3��y ��Ɏ����H8�o�0�z~�sPD��X��Q��@�d�z��k�y "���&i�SOI��~S�!�Ĺ"z��%f��ʆ3ߞK�J�,o���x�Z!���W�NkpyR�G[���ѣ^<�gq)�T87`\��/�B�rk^�g��[.2h�g�;ҙ2��a57�9^�Ž�[I�?��K"^��@�}�mx�R��&���6�=�GP]�j=�߼H._�-m��)�H6Q!�I��6��
'���n�08�U@����9�pd�5�(�н�K��gr����y_jҁ��Vh�z����#����Q G6�u�
��*�2���pu�'Y�W�c�~qO�)�1	b�+���U�|�qK���������8?㘰�,�S��O[{���]k�A%�*��6�Y���-�M��Z�C<��~	 �$��4B}@��&�	O���������������L����գh���J�^�;g.��W�3l�=3�G1Q�A�f�<AIooͥ������	1��^׻�����Y��m��?z�6����0��V|~ךa��J0����Wr|�/�zv\$�S�H�[��N�R�G7r�v�9�,�*�ؕ���Qh���,�£��n�8/ⱖs$�My^��P΅7^���Z�	���-���G��Z?;�m� sA�E��L�S�~�C�V^��YW-U|���Z��}�2t��f�] ���n"�k(�K����r�\JTa�f��~�����3ak' M:��"�GB��Ud?$Xt���p�J�y����l]&�h��E� �L\���<y^�:������/�������֥Rq���d�/n�s�	Hg��j�g�&��;�?��3r�}���թ�9������YU���_��:m�F���
j���"�e��A0��^Е���g�P;,����tn�]�v�cH�M=�^�]��ΩaydI�2ݰ�!Hk�R:_6Sx��b�/�-ZE�}��EJ�fz*��Q������y�Ua9�M w�?Yy�����=�k�aĂ�~��]	���t1ʩs��oC��#��L��A/�� �p)����~��D�ߣT��k�R�?�{m�'Ѱ�dR~ ��I{��YӜI˂��^�J��,��W����X����oG���/P�,;��*�k8�N&Z��.���#3-F��	Y�/���	&UEpok�U��s(��{RY��f"����&��?�������7hs�N�n5~�ɋ��  �%�|r���#�s�.��+�h��\D���ں�-�L�}&�
�Vt/c�#���J����e☘f@A�������U� `rɳ%�h� _��n�GIt�G#Ì�~�-&�
�ѯ2A�g[ RHN�"����P�wFL/�h6�>��ޭ�W� p
��0�Vv����c;�
�K�Q����<O�s�F>��@k-��Y����&��ڌ����͂��Ed���ؤ�8:�|�
3{je�����*!u4��mg!S?��a�uZR��S<�=���֘w����i'�nԛY��	���8�|
�E
[U�qT��yċ-�kyx�ړ���� T��)U�RX�;e
��e�tMJO��?U�IS����;��G\��~��8�7��;��?��L�']<� �s��I�tl�g9�����%��^B�mE��S���2e��J����b��<]S�wz��
\�ߏ�*c�r�l������o���?��P����Ă��-��W��nS��k��t$����\�J䓋�Ӏ����#�}���Gs�P*lt=f�������������&B���$41���jh?l��;��$%���=�W����ʴb��#\���^�
�d�#�2������j�C;�S<��ǽ�q���H��=y�~rTة�M�`Q�[��j�iۦ�T�\PG����f���tgU�:Z���Zțcd��M��:�h��X�����Q���E�;c�8�$���_A}����]�'`~~V���۲����wR�H,�2~r�����AY�h/����zeZ�G%^/����G��>��]��Z^k�$j�L�����G��B��r_uf��Ӊ�0�E�0Gto�ㆃ��^�0/=2�ʺ�����C�E�*	]t�G�o���p���o����C���o�$#�R��z=�U{^��{�Sr�DRo��� W�g�K�<��*���J,����R��;��h�ڃ�q���
���8��&�B��?"���<���p���b@�#FUE>��������&���G�y`�W�	�r�$�wSv�q+/ב�4���M4p�-���p��`�8�>�k�����>�q��_�e@E�z�%n�?n�6l"�L A�\�(M�P��Kb������h�/*�I!b���Oe�l��I2}�d��G/{��=K2a���f7ߴ��ހ��'6D����B'�o�$s�?��`��&��Rw�����n�`;ӧ᫏r�V8.�r�8�He��Y��^�4:A
 ���9�/�R*�A�_�z%����]b,>|x�W���KTb��AS����d8P�`8�Q]q�f�Ӽ�k&�[h�Œ./�k�os~�����¾Қ_Ԩ�>��	H�n:}ksݟ����=g<y�O����Ia�W.|�gB|{�o�Rb2��%�Q���9�L
��=���.���;��T���ݥvp1���C&�W$�  �o^q�!1�����@;��]���Ɗ�S�a��d�$����%��7�)d2�v�~�C�ݿ$J�&�"�,�sʬ�|aK�+U�vD�<ԾHÍ�
��*�PڋJ�6��bU}�<��w(��/�ժ�&[#_X�2��zN�{S�|�p��a��pu­/��8����z(Qd��Mb��n�]�ӫ�f���)��q�?�?�r����,�b�,S��aw����X|(_��m��'� qee!��n�X Q�h��`��3|�ɷB�&4����2hr��7��Xr~�"e�����5s%$�'�c��DඩT�!�����r{�[�v�Ѥ��
w#GM�Q�H�kH�L`j.,9������5=�Kn��k�OC�G�������PT�c�(��g=O���og�[w�
���Գ�� �D�JJ�!O��n,UE+�},�k��y[z�i%'r�[�n� O]��e�/�ğ�p�d8�P/;m">~��hz>���PQ�w��D`:��,/�����<�M�Aќ����G�Ч,{I�J+e�s��%C���wz
�EiX@+G�+c\6c�j���J��n�c0���GI>������ bTÇ,p�{���tn�N�A��LW�c��x�Xh�P%�%�����{�y�R��)���7��ՙ֣�F@A�]}Cmo�#>���."][+�������I��JLkC���o�4�h-go�K�:���Ɂ/��Y�㥄�yv#��2�w��g��8�S�@��d�ұ�t�C��9I��-��&]�6s�i��:����R/'�a�x��$3ІI��!O�i?�:��	J��n������IH4�����1Q�28`���@��5��*�]d�ak�5��M&==g�GS9Q��A��-�	F��5�X��7�y�a�����-7U~|���ez�N�^o@�kE(6&����fL����������0�[/��$�A��9<�`@���Sc�7&1�Oik8��3����`v�3'j*���!��Ɨ�(E�l%���mk�<_��<���7�a��Ȭ\g���:�\�g"F9m^���çN�@�����k�D;3����vkp�&�*��֥;W��а~{4�F�5�Zr��E�(d�����+���1A�9���n^�%F��m%�IQ����Η-�2������Q>�9`;F��l�ӘN�?� ��"�����	�3���ux��\}*e�9n  ��OG�����wA�Y��nO�B�^S�1�qȂX�/#��Vk��p�T�l5�&	�	n�p�m]��b� 3u��{�[���k�fX�\��?�`�E�wO{Q*A&*@�D@�7�R��IGF~/fF�Ҥ/z��N�����p� ۭ�Zy�Arɮ�3�ڥ>�b����q�H&�3xe��;�^�0�-Y	��jl��Z���.�:c�?+]�"С��7��&Q�@|�I2ȱ<<CHƧx=s=Rs�b3n�=5�mJG-�3d]�f��Ja3|���"�-�jǩ�G�4)N���P\.��Nq�VH�ݎ[���*%N�4L����*�ARA�>>.V�Ք�'Tq��>�,sG~�N 1��y�o��:Nw�vi�Y7T�����2�\�L��m�U�@������� D��9��)����.Q�i���]�q�aU��T�@{6��=#�d^Xt���A�%P ��Mi����;Զ�W��鏊vH�?�C$u�}�U2���pd��*����/1���8�e�5��Ȇ=����G9`��_-H���O�0���m���%�S���j��&��ј���������_a�	=�ie�0���!��,��y�)+��.2N�2��z-�Pؗ��;J(*:%gdF*�(���h�5] m���rj�K�{��Q2<6���@AO��n1�s��KoO���_��RJ#B��+\d�Uݩ�[��{��n��j�p�ZGqA#g��㒊F��S�.5{8i�}̹�s^�e���F|�!��T$9q��Ko�,D`�S�PaN*�M<'����nZ��������O\4~Y�Sx�n`�=�I��T�⯷���K<���r�A$�ý�Yރ���%F�T�ez��/!��f�K&����R5�N�	����B�V6�'E���-������V�
��@#���	-��xx�����i��(;~0����A��:2�)Y}+B�^��qf��/�M���s�RkO�%�$�8��2�u�7,J���}����)�k�vN���Z�V	Y�%�ϛ��d��/��`(��L'�I�T���*�RJ`���#�� h|7�˟�|�-ev4T0 �ٝs7I9�%1�������ݨ}x�-Щ�i����R���R�@�25���#�r�ՠ�~4a2psÂQ��!oY��H��;Z6u�p�Z�iڷ�?����6���A���a�$bl��)O�� ��a���7�Y����Di��Pų��ʗgtt�M��;���?�#Ďg�T��f�ۇ\	�H
�	4��/SŚ~���m�Ҫz�?-���ޝ�~@a���lʐ+���Y"<�>X��\3s�BF?�=�Lr1 ipp�d�,�'�t��Uf��E��$L=Qǀu5�zf�
-��5�Riэ��sC�<��Gc.T�fjep���^�-]t�'s����X�̇�I}e�a��� '�u�:wԬ�,d���z�/�	T1�+�O���=�Ǆ����D�
e�L��(F'�W����}ߗxX2�z�{�3�tN%���{k����G�VA<}d�����Y�ք���n,����I�=�Z�j�����o����J��C�Hxt�w��{!	Ck�u��:�Ig���fʡ	�-����@T��t��"��S4Ne��X6����:<���@�$��E�%Z������t��dHh���h1B��!U�������r@�]�^��qZ�i {!j_�Ѝ1���@$ Jm�
e�
�_�������eP����XFz	[Q�eԯ_��1Z-�Ifg4* c�Ͷ����"�����g�r��.����p�Q6q>��>G��%��>V07�xO�����{���;ϳ��afyс�$LX�ּ7�&�O���ҏ�u��9�O�F���:bWu�[���	LD!u4���~ؖ��V�
҉�ɋ/�Ϙ��T_�{��?i�K̟�9iG��&�CV	v��0 
w�PV}�y�+���24F�y\/������_H��#�g�����Q��9���tGV�,m�Ӌ{G�J��x�VOEa�˧;����}��ۗ�=ө��]<7
y�8���@�5���!����#ILr��Q�����l��]��	�Y=�^��JTj� ������ݵejTj�ʐ�}�e#B�#��x�C������Bj�C���P߬Wt(e������:AK�:\�a�ii*ְ��I�$zE ��_e���k;��Z���د��gm(�<���0��Y���ba,�Sq�H�F%�$��vǢ�=��6����u9�Ī=��{ܗ^�M��lՇrs�����#͇A8u��~���4�K_�x����Y4��*K�/��z����[H����qxAb�(*T3P��ü��=U�R��A�f!����Z³&G����Kv�=
�L):�2���#�!2�������Ulr��NTsAD�)�O�/�^�G"&U�%�3]o�	X�E ^�Y�2R�X��eq9�Ŝ��V��T*��A�����[�v�`3�-�!��n�^����:k�<4#v�\t��3�r	�>���D���o2�n�d�*�����ó~g.�v1N)�Ɩ����
� �-����p��u%B��.{1Xo{�371�j�����k퍃�
���D8����!0J�_;��ӊ5���lo�k���j��A�����OpA���f3�3Vʢ+w�أ��|���X}���
�C�!�ŧ7�O��z���h�l��ԠQ�>�(U}���Z^�U�$�ì���2�g�ڥ��ⵧ�?���3k�м��Ӿ*��7SY��O����G��Y����"�o�8]̮,e��t7�j����G��� t���^0!)��X}��3(foS���H5�<�B��k0�D"�e����7Ա�S��d(}�T*g��	�ʇ�{��'��ZNŰ��#�}��
�ცA��	ʞ�ْ]���\3�����jGqY㋈�`��YFq(�Ue��P�ִpz�,�Q�mB<y-X]��6�:ש�lT�����bP��-F��k��ˡ��c�,1�)ťx�WK*��E�
��܈5٬�YC5�3���
�T>������I������kx�$�~�{�$�	>�� �n��e����b�#���P��cI����JM0�̃�N�G��>ئg���[ɯ�^N4���ō�����+�8���κs�ۼ�m��2h�^�Du����Ğ�R"�cE 7�S 啔�q{I�����G���4R�D�.�'M�UI+Z\��&,�������!ﺮ�H�7������~c��;tQ�Z��Tt�Ʋ+%�#tg�#m����Qj��G�8&����bP]0�.C�.�$ ��À�|3�bq�}����hyh5�;�`�.�����"�+�	 �_�� }:�C��5��a��B캯���1LQe�9}�4��KUI����*'�`1�Pd(7���FR&i��9��vԓ�}"�n�MÈu�Wg���?��t��8p���E؉Q��q�0s����k�Ƙ̽U3N�K��/E�j��H�\�q���?g��\X-~�E�z.ɪo��4k�x[\�l��b�ɥa�2Kx.�Xhj�)i���tH�yũ�:��p��LM��Jq��.��t��#-����7@\<U,�%�C�,9!sWy��Ҡq������6b����r�_���]~yx�f����Z�(�M]u}���ܪNG��j4�3�S;q���p
ݭ��z��#:Ү�"NI	�?�53R�"�����n�e��,}�˦���q�·����ͳcE�c�렪�<\�I��J����Ϥ�И��s���3jp�.��u,O���l�3��NL7	8�U
��������=�1�p&,
Ĩ�/&b8�¨m�Q���Z��D��{yKo@��'Q�q��i���{���دGTΔ��LY�8[�jS��3��VO��I�$m2x�����h�!̪��w�(�0�.�s�*��M�C�s�>��F��;ݵ���	d�H��*�� ��,?6~�L�A���1e5,���f�</�Rz��z9��>�&k;���R�u#�^�j��9��q����9UO�Z+��X��奕 #�#0R��L"��[��4��f�[�Ǯv�W�i����$�}�(�:�Ӗ���("�LZ�QL�����_��r�������r��R��ض��νnv!��?�{uh�sR�v�_˟TseCs���	�� ��{�>���V�;��⋸���mTF��p�Hͬ�d)�E��˖�d#�1�/8 �|�|�eFU�-��0���x�7-�l*�`��l��hL:;��O�Z-1j�?b����4r��+�L������L���q͢=��<�c"Vf�������r��w��5����f'Ӂzo�i�>#�
�x*���h�+